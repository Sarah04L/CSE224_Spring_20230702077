VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cpu_lab6
  CLASS BLOCK ;
  FOREIGN cpu_lab6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 100.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 11.020 10.640 12.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.020 10.640 32.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.020 10.640 52.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.020 10.640 72.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.020 10.640 92.620 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 16.380 94.540 17.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 36.380 94.540 37.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 56.380 94.540 57.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 76.380 94.540 77.980 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 7.720 10.640 9.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 27.720 10.640 29.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.720 10.640 49.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 67.720 10.640 69.320 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 87.720 10.640 89.320 87.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 13.080 94.540 14.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 33.080 94.540 34.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 53.080 94.540 54.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 73.080 94.540 74.680 ;
    END
  END VPWR
  PIN an[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END an[0]
  PIN an[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END an[1]
  PIN an[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END an[2]
  PIN an[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END an[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END clk
  PIN control
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END control
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END reset
  PIN seg[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END seg[0]
  PIN seg[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 51.040 100.000 51.640 ;
    END
  END seg[1]
  PIN seg[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END seg[2]
  PIN seg[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 96.000 48.670 100.000 ;
    END
  END seg[3]
  PIN seg[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 96.000 51.890 100.000 ;
    END
  END seg[4]
  PIN seg[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END seg[5]
  PIN seg[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END seg[6]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 94.490 87.125 ;
      LAYER li1 ;
        RECT 5.520 10.795 94.300 87.125 ;
      LAYER met1 ;
        RECT 4.210 10.640 94.300 87.280 ;
      LAYER met2 ;
        RECT 4.230 95.720 48.110 96.000 ;
        RECT 48.950 95.720 51.330 96.000 ;
        RECT 52.170 95.720 92.830 96.000 ;
        RECT 4.230 4.280 92.830 95.720 ;
        RECT 4.230 4.000 6.250 4.280 ;
        RECT 7.090 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 92.830 4.280 ;
      LAYER met3 ;
        RECT 3.990 58.840 96.000 87.205 ;
        RECT 4.400 57.440 96.000 58.840 ;
        RECT 3.990 55.440 96.000 57.440 ;
        RECT 4.400 54.040 96.000 55.440 ;
        RECT 3.990 52.040 96.000 54.040 ;
        RECT 4.400 50.640 95.600 52.040 ;
        RECT 3.990 48.640 96.000 50.640 ;
        RECT 4.400 47.240 96.000 48.640 ;
        RECT 3.990 45.240 96.000 47.240 ;
        RECT 4.400 43.840 96.000 45.240 ;
        RECT 3.990 41.840 96.000 43.840 ;
        RECT 4.400 40.440 96.000 41.840 ;
        RECT 3.990 10.715 96.000 40.440 ;
  END
END cpu_lab6
END LIBRARY

