module myBasic_ALU (A,
    B,
    opcode,
    out);
 input [7:0] A;
 input [7:0] B;
 input [2:0] opcode;
 output [8:0] out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;

 sky130_fd_sc_hd__clkbuf_2 _170_ (.A(net4),
    .X(_100_));
 sky130_fd_sc_hd__or2_1 _171_ (.A(net17),
    .B(net18),
    .X(_101_));
 sky130_fd_sc_hd__nor2_2 _172_ (.A(net19),
    .B(_101_),
    .Y(_102_));
 sky130_fd_sc_hd__buf_2 _173_ (.A(_102_),
    .X(_103_));
 sky130_fd_sc_hd__buf_2 _174_ (.A(net3),
    .X(_104_));
 sky130_fd_sc_hd__buf_2 _175_ (.A(net11),
    .X(_105_));
 sky130_fd_sc_hd__nand3b_4 _176_ (.A_N(net17),
    .B(net18),
    .C(net19),
    .Y(_106_));
 sky130_fd_sc_hd__or2_1 _177_ (.A(net10),
    .B(net9),
    .X(_107_));
 sky130_fd_sc_hd__nand2_1 _178_ (.A(net29),
    .B(_107_),
    .Y(_108_));
 sky130_fd_sc_hd__xor2_1 _179_ (.A(_105_),
    .B(_108_),
    .X(_109_));
 sky130_fd_sc_hd__and2_1 _180_ (.A(_104_),
    .B(_109_),
    .X(_110_));
 sky130_fd_sc_hd__buf_2 _181_ (.A(net10),
    .X(_111_));
 sky130_fd_sc_hd__buf_2 _182_ (.A(net9),
    .X(_112_));
 sky130_fd_sc_hd__and3_1 _183_ (.A(_111_),
    .B(_112_),
    .C(_106_),
    .X(_113_));
 sky130_fd_sc_hd__a21oi_1 _184_ (.A1(_112_),
    .A2(_106_),
    .B1(_111_),
    .Y(_114_));
 sky130_fd_sc_hd__or3_4 _185_ (.A(net2),
    .B(_113_),
    .C(_114_),
    .X(_115_));
 sky130_fd_sc_hd__inv_2 _186_ (.A(net1),
    .Y(_116_));
 sky130_fd_sc_hd__nand2_1 _187_ (.A(_116_),
    .B(_112_),
    .Y(_117_));
 sky130_fd_sc_hd__o21a_1 _188_ (.A1(_113_),
    .A2(_114_),
    .B1(net2),
    .X(_118_));
 sky130_fd_sc_hd__a21o_1 _189_ (.A1(_117_),
    .A2(_115_),
    .B1(_118_),
    .X(_119_));
 sky130_fd_sc_hd__xor2_1 _190_ (.A(_104_),
    .B(_109_),
    .X(_120_));
 sky130_fd_sc_hd__and2_4 _191_ (.A(_119_),
    .B(_120_),
    .X(_121_));
 sky130_fd_sc_hd__o21a_1 _192_ (.A1(net11),
    .A2(_107_),
    .B1(net29),
    .X(_122_));
 sky130_fd_sc_hd__xnor2_1 _193_ (.A(net12),
    .B(_122_),
    .Y(_123_));
 sky130_fd_sc_hd__and2_1 _194_ (.A(_100_),
    .B(_123_),
    .X(_124_));
 sky130_fd_sc_hd__or2_1 _195_ (.A(_100_),
    .B(_123_),
    .X(_125_));
 sky130_fd_sc_hd__and2b_1 _196_ (.A_N(_124_),
    .B(_125_),
    .X(_126_));
 sky130_fd_sc_hd__o21ai_1 _197_ (.A1(_110_),
    .A2(_121_),
    .B1(_126_),
    .Y(_127_));
 sky130_fd_sc_hd__nand2_1 _198_ (.A(net17),
    .B(net18),
    .Y(_128_));
 sky130_fd_sc_hd__and3_2 _199_ (.A(net19),
    .B(_101_),
    .C(_128_),
    .X(_129_));
 sky130_fd_sc_hd__o31a_1 _200_ (.A1(_126_),
    .A2(_110_),
    .A3(_121_),
    .B1(_129_),
    .X(_130_));
 sky130_fd_sc_hd__nand2_1 _201_ (.A(_105_),
    .B(net1),
    .Y(_131_));
 sky130_fd_sc_hd__and2_1 _202_ (.A(net2),
    .B(_112_),
    .X(_132_));
 sky130_fd_sc_hd__and2_1 _203_ (.A(net10),
    .B(net3),
    .X(_133_));
 sky130_fd_sc_hd__a22o_1 _204_ (.A1(net10),
    .A2(net2),
    .B1(net3),
    .B2(_112_),
    .X(_134_));
 sky130_fd_sc_hd__a21bo_1 _205_ (.A1(_132_),
    .A2(_133_),
    .B1_N(_134_),
    .X(_135_));
 sky130_fd_sc_hd__xor2_1 _206_ (.A(_131_),
    .B(_135_),
    .X(_136_));
 sky130_fd_sc_hd__and3_1 _207_ (.A(_111_),
    .B(net1),
    .C(_132_),
    .X(_137_));
 sky130_fd_sc_hd__and2_1 _208_ (.A(_136_),
    .B(_137_),
    .X(_138_));
 sky130_fd_sc_hd__buf_2 _209_ (.A(net12),
    .X(_139_));
 sky130_fd_sc_hd__nand2_1 _210_ (.A(_139_),
    .B(net1),
    .Y(_140_));
 sky130_fd_sc_hd__o2bb2a_1 _211_ (.A1_N(_132_),
    .A2_N(_133_),
    .B1(_135_),
    .B2(_131_),
    .X(_141_));
 sky130_fd_sc_hd__nand2_1 _212_ (.A(_105_),
    .B(net2),
    .Y(_142_));
 sky130_fd_sc_hd__nand4_1 _213_ (.A(net4),
    .B(_111_),
    .C(net3),
    .D(_112_),
    .Y(_143_));
 sky130_fd_sc_hd__a22o_1 _214_ (.A1(_111_),
    .A2(net3),
    .B1(_112_),
    .B2(net4),
    .X(_144_));
 sky130_fd_sc_hd__nand2_1 _215_ (.A(_143_),
    .B(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__xor2_1 _216_ (.A(_142_),
    .B(_145_),
    .X(_146_));
 sky130_fd_sc_hd__xnor2_1 _217_ (.A(_141_),
    .B(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__xnor2_1 _218_ (.A(_140_),
    .B(_147_),
    .Y(_148_));
 sky130_fd_sc_hd__and2_1 _219_ (.A(_138_),
    .B(_148_),
    .X(_149_));
 sky130_fd_sc_hd__inv_2 _220_ (.A(net19),
    .Y(_150_));
 sky130_fd_sc_hd__nor2_2 _221_ (.A(_150_),
    .B(_101_),
    .Y(_151_));
 sky130_fd_sc_hd__o21ai_1 _222_ (.A1(_138_),
    .A2(_148_),
    .B1(_151_),
    .Y(_152_));
 sky130_fd_sc_hd__nor2_2 _223_ (.A(net19),
    .B(_128_),
    .Y(_153_));
 sky130_fd_sc_hd__nand2_1 _224_ (.A(net17),
    .B(_150_),
    .Y(_154_));
 sky130_fd_sc_hd__nor2_2 _225_ (.A(net18),
    .B(_154_),
    .Y(_155_));
 sky130_fd_sc_hd__or3b_1 _226_ (.A(net17),
    .B(net19),
    .C_N(net18),
    .X(_156_));
 sky130_fd_sc_hd__clkbuf_2 _227_ (.A(_156_),
    .X(_157_));
 sky130_fd_sc_hd__a21oi_1 _228_ (.A1(_100_),
    .A2(_139_),
    .B1(_157_),
    .Y(_158_));
 sky130_fd_sc_hd__o22a_1 _229_ (.A1(_100_),
    .A2(_139_),
    .B1(_155_),
    .B2(_158_),
    .X(_159_));
 sky130_fd_sc_hd__a311o_1 _230_ (.A1(_100_),
    .A2(_139_),
    .A3(_153_),
    .B1(_159_),
    .C1(_102_),
    .X(_160_));
 sky130_fd_sc_hd__o21bai_1 _231_ (.A1(_149_),
    .A2(_152_),
    .B1_N(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__a21oi_1 _232_ (.A1(_127_),
    .A2(_130_),
    .B1(_161_),
    .Y(_162_));
 sky130_fd_sc_hd__a21oi_1 _233_ (.A1(_100_),
    .A2(_103_),
    .B1(_162_),
    .Y(net23));
 sky130_fd_sc_hd__nand2_1 _234_ (.A(net12),
    .B(net2),
    .Y(_163_));
 sky130_fd_sc_hd__a22oi_1 _235_ (.A1(net4),
    .A2(_111_),
    .B1(_104_),
    .B2(_105_),
    .Y(_164_));
 sky130_fd_sc_hd__and3_1 _236_ (.A(net4),
    .B(net11),
    .C(_133_),
    .X(_165_));
 sky130_fd_sc_hd__or2_1 _237_ (.A(_164_),
    .B(_165_),
    .X(_166_));
 sky130_fd_sc_hd__o21ai_1 _238_ (.A1(_142_),
    .A2(_145_),
    .B1(_143_),
    .Y(_167_));
 sky130_fd_sc_hd__xnor2_1 _239_ (.A(_166_),
    .B(_167_),
    .Y(_168_));
 sky130_fd_sc_hd__xnor2_1 _240_ (.A(_163_),
    .B(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__and2b_1 _241_ (.A_N(_141_),
    .B(_146_),
    .X(_000_));
 sky130_fd_sc_hd__a31o_1 _242_ (.A1(_139_),
    .A2(net1),
    .A3(_147_),
    .B1(_000_),
    .X(_001_));
 sky130_fd_sc_hd__xor2_1 _243_ (.A(_169_),
    .B(_001_),
    .X(_002_));
 sky130_fd_sc_hd__xor2_1 _244_ (.A(_149_),
    .B(_002_),
    .X(_003_));
 sky130_fd_sc_hd__o31a_1 _245_ (.A1(net12),
    .A2(_105_),
    .A3(_107_),
    .B1(net30),
    .X(_004_));
 sky130_fd_sc_hd__xnor2_1 _246_ (.A(_004_),
    .B(net13),
    .Y(_005_));
 sky130_fd_sc_hd__and2_4 _247_ (.A(_005_),
    .B(net5),
    .X(_006_));
 sky130_fd_sc_hd__nor2_1 _248_ (.A(net5),
    .B(_005_),
    .Y(_007_));
 sky130_fd_sc_hd__nor2_1 _249_ (.A(_006_),
    .B(_007_),
    .Y(_008_));
 sky130_fd_sc_hd__or2_1 _250_ (.A(_124_),
    .B(_110_),
    .X(_009_));
 sky130_fd_sc_hd__o21a_1 _251_ (.A1(_121_),
    .A2(_009_),
    .B1(_125_),
    .X(_010_));
 sky130_fd_sc_hd__or2_1 _252_ (.A(_008_),
    .B(_010_),
    .X(_011_));
 sky130_fd_sc_hd__o211a_4 _253_ (.A1(_121_),
    .A2(_009_),
    .B1(_008_),
    .C1(_125_),
    .X(_012_));
 sky130_fd_sc_hd__and2b_1 _254_ (.A_N(_012_),
    .B(_129_),
    .X(_013_));
 sky130_fd_sc_hd__a21oi_1 _255_ (.A1(net5),
    .A2(net13),
    .B1(_157_),
    .Y(_014_));
 sky130_fd_sc_hd__o22a_1 _256_ (.A1(net5),
    .A2(net13),
    .B1(_155_),
    .B2(_014_),
    .X(_015_));
 sky130_fd_sc_hd__a311o_1 _257_ (.A1(net5),
    .A2(net13),
    .A3(_153_),
    .B1(_015_),
    .C1(_102_),
    .X(_016_));
 sky130_fd_sc_hd__a21o_1 _258_ (.A1(_011_),
    .A2(_013_),
    .B1(_016_),
    .X(_017_));
 sky130_fd_sc_hd__a21oi_1 _259_ (.A1(_151_),
    .A2(_003_),
    .B1(_017_),
    .Y(_018_));
 sky130_fd_sc_hd__a21oi_1 _260_ (.A1(net5),
    .A2(_103_),
    .B1(_018_),
    .Y(net24));
 sky130_fd_sc_hd__o41a_1 _261_ (.A1(net12),
    .A2(net13),
    .A3(net11),
    .A4(_107_),
    .B1(net30),
    .X(_019_));
 sky130_fd_sc_hd__xor2_1 _262_ (.A(net14),
    .B(_019_),
    .X(_020_));
 sky130_fd_sc_hd__or2b_2 _263_ (.A(net6),
    .B_N(_020_),
    .X(_021_));
 sky130_fd_sc_hd__inv_2 _264_ (.A(_021_),
    .Y(_022_));
 sky130_fd_sc_hd__and2b_1 _265_ (.A_N(_020_),
    .B(net6),
    .X(_023_));
 sky130_fd_sc_hd__nor2_1 _266_ (.A(_022_),
    .B(_023_),
    .Y(_024_));
 sky130_fd_sc_hd__o21ai_1 _267_ (.A1(_006_),
    .A2(_012_),
    .B1(_024_),
    .Y(_025_));
 sky130_fd_sc_hd__o31a_1 _268_ (.A1(_006_),
    .A2(_012_),
    .A3(_024_),
    .B1(_129_),
    .X(_026_));
 sky130_fd_sc_hd__and2_1 _269_ (.A(_025_),
    .B(_026_),
    .X(_027_));
 sky130_fd_sc_hd__or2b_1 _270_ (.A(_166_),
    .B_N(_167_),
    .X(_028_));
 sky130_fd_sc_hd__or2b_1 _271_ (.A(_163_),
    .B_N(_168_),
    .X(_029_));
 sky130_fd_sc_hd__and3b_1 _272_ (.A_N(_133_),
    .B(_105_),
    .C(_100_),
    .X(_030_));
 sky130_fd_sc_hd__nand2_1 _273_ (.A(_139_),
    .B(_104_),
    .Y(_031_));
 sky130_fd_sc_hd__xor2_1 _274_ (.A(_030_),
    .B(_031_),
    .X(_032_));
 sky130_fd_sc_hd__and3_1 _275_ (.A(_028_),
    .B(_029_),
    .C(_032_),
    .X(_033_));
 sky130_fd_sc_hd__a21oi_1 _276_ (.A1(_028_),
    .A2(_029_),
    .B1(_032_),
    .Y(_034_));
 sky130_fd_sc_hd__nor2_1 _277_ (.A(_033_),
    .B(_034_),
    .Y(_035_));
 sky130_fd_sc_hd__nand2_1 _278_ (.A(_169_),
    .B(_001_),
    .Y(_036_));
 sky130_fd_sc_hd__a21boi_1 _279_ (.A1(_149_),
    .A2(_002_),
    .B1_N(_036_),
    .Y(_037_));
 sky130_fd_sc_hd__xnor2_1 _280_ (.A(_035_),
    .B(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__a21oi_1 _281_ (.A1(net6),
    .A2(net14),
    .B1(_157_),
    .Y(_039_));
 sky130_fd_sc_hd__o22a_1 _282_ (.A1(net6),
    .A2(net14),
    .B1(_155_),
    .B2(_039_),
    .X(_040_));
 sky130_fd_sc_hd__a31o_1 _283_ (.A1(net6),
    .A2(net14),
    .A3(_153_),
    .B1(_040_),
    .X(_041_));
 sky130_fd_sc_hd__a211o_1 _284_ (.A1(_151_),
    .A2(_038_),
    .B1(_041_),
    .C1(_103_),
    .X(_042_));
 sky130_fd_sc_hd__o2bb2a_1 _285_ (.A1_N(net6),
    .A2_N(_103_),
    .B1(_027_),
    .B2(_042_),
    .X(net25));
 sky130_fd_sc_hd__a21o_1 _286_ (.A1(net14),
    .A2(net31),
    .B1(_019_),
    .X(_043_));
 sky130_fd_sc_hd__xnor2_1 _287_ (.A(net15),
    .B(_043_),
    .Y(_044_));
 sky130_fd_sc_hd__nand2_1 _288_ (.A(net7),
    .B(_044_),
    .Y(_045_));
 sky130_fd_sc_hd__or2_1 _289_ (.A(net7),
    .B(_044_),
    .X(_046_));
 sky130_fd_sc_hd__and2_4 _290_ (.A(_045_),
    .B(_046_),
    .X(_047_));
 sky130_fd_sc_hd__o31a_1 _291_ (.A1(_006_),
    .A2(_012_),
    .A3(_023_),
    .B1(_021_),
    .X(_048_));
 sky130_fd_sc_hd__or2_1 _292_ (.A(_047_),
    .B(_048_),
    .X(_049_));
 sky130_fd_sc_hd__o311ai_4 _293_ (.A1(_006_),
    .A2(_023_),
    .A3(_012_),
    .B1(_047_),
    .C1(_021_),
    .Y(_050_));
 sky130_fd_sc_hd__and3_1 _294_ (.A(_129_),
    .B(_049_),
    .C(_050_),
    .X(_051_));
 sky130_fd_sc_hd__a31o_1 _295_ (.A1(_139_),
    .A2(_104_),
    .A3(_030_),
    .B1(_165_),
    .X(_052_));
 sky130_fd_sc_hd__a21oi_1 _296_ (.A1(_100_),
    .A2(_139_),
    .B1(_052_),
    .Y(_053_));
 sky130_fd_sc_hd__a41o_1 _297_ (.A1(_100_),
    .A2(_139_),
    .A3(_105_),
    .A4(_104_),
    .B1(_053_),
    .X(_054_));
 sky130_fd_sc_hd__o21ba_1 _298_ (.A1(_036_),
    .A2(_033_),
    .B1_N(_034_),
    .X(_055_));
 sky130_fd_sc_hd__xor2_1 _299_ (.A(_054_),
    .B(_055_),
    .X(_056_));
 sky130_fd_sc_hd__a21oi_1 _300_ (.A1(net7),
    .A2(net15),
    .B1(_157_),
    .Y(_057_));
 sky130_fd_sc_hd__o22a_1 _301_ (.A1(net7),
    .A2(net15),
    .B1(_155_),
    .B2(_057_),
    .X(_058_));
 sky130_fd_sc_hd__a31o_1 _302_ (.A1(net7),
    .A2(net15),
    .A3(_153_),
    .B1(_058_),
    .X(_059_));
 sky130_fd_sc_hd__a211o_1 _303_ (.A1(_151_),
    .A2(_056_),
    .B1(_059_),
    .C1(_102_),
    .X(_060_));
 sky130_fd_sc_hd__o2bb2a_1 _304_ (.A1_N(net7),
    .A2_N(_103_),
    .B1(_051_),
    .B2(_060_),
    .X(net26));
 sky130_fd_sc_hd__o21a_1 _305_ (.A1(net15),
    .A2(_043_),
    .B1(net31),
    .X(_061_));
 sky130_fd_sc_hd__xnor2_1 _306_ (.A(net16),
    .B(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__xor2_1 _307_ (.A(net8),
    .B(_062_),
    .X(_063_));
 sky130_fd_sc_hd__inv_2 _308_ (.A(_063_),
    .Y(_064_));
 sky130_fd_sc_hd__nand3_1 _309_ (.A(_045_),
    .B(_050_),
    .C(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__a21o_1 _310_ (.A1(_045_),
    .A2(_050_),
    .B1(_064_),
    .X(_066_));
 sky130_fd_sc_hd__and3_1 _311_ (.A(_129_),
    .B(_065_),
    .C(_066_),
    .X(_067_));
 sky130_fd_sc_hd__nand3_1 _312_ (.A(_100_),
    .B(_139_),
    .C(_052_),
    .Y(_068_));
 sky130_fd_sc_hd__o21ai_1 _313_ (.A1(_053_),
    .A2(_055_),
    .B1(_068_),
    .Y(_069_));
 sky130_fd_sc_hd__a21oi_1 _314_ (.A1(net8),
    .A2(net16),
    .B1(_157_),
    .Y(_070_));
 sky130_fd_sc_hd__o22a_1 _315_ (.A1(net8),
    .A2(net16),
    .B1(_155_),
    .B2(_070_),
    .X(_071_));
 sky130_fd_sc_hd__a31o_1 _316_ (.A1(net8),
    .A2(net16),
    .A3(_153_),
    .B1(_071_),
    .X(_072_));
 sky130_fd_sc_hd__a211o_1 _317_ (.A1(_151_),
    .A2(_069_),
    .B1(_072_),
    .C1(_102_),
    .X(_073_));
 sky130_fd_sc_hd__o2bb2a_1 _318_ (.A1_N(net8),
    .A2_N(_103_),
    .B1(_067_),
    .B2(_073_),
    .X(net27));
 sky130_fd_sc_hd__and3b_1 _319_ (.A_N(net17),
    .B(net18),
    .C(net19),
    .X(_074_));
 sky130_fd_sc_hd__nor2_1 _320_ (.A(net16),
    .B(_061_),
    .Y(_075_));
 sky130_fd_sc_hd__nand2_1 _321_ (.A(net8),
    .B(_062_),
    .Y(_076_));
 sky130_fd_sc_hd__a2bb2o_1 _322_ (.A1_N(_074_),
    .A2_N(_075_),
    .B1(_076_),
    .B2(_066_),
    .X(_077_));
 sky130_fd_sc_hd__or4bb_1 _323_ (.A(_074_),
    .B(_075_),
    .C_N(_076_),
    .D_N(_066_),
    .X(_078_));
 sky130_fd_sc_hd__a31o_1 _324_ (.A1(_129_),
    .A2(_077_),
    .A3(_078_),
    .B1(_103_),
    .X(net28));
 sky130_fd_sc_hd__or2_1 _325_ (.A(net1),
    .B(_112_),
    .X(_079_));
 sky130_fd_sc_hd__nand3_1 _326_ (.A(net1),
    .B(_112_),
    .C(_154_),
    .Y(_080_));
 sky130_fd_sc_hd__o211a_1 _327_ (.A1(_151_),
    .A2(_153_),
    .B1(net1),
    .C1(_112_),
    .X(_081_));
 sky130_fd_sc_hd__a31o_1 _328_ (.A1(_101_),
    .A2(_128_),
    .A3(_080_),
    .B1(_081_),
    .X(_082_));
 sky130_fd_sc_hd__a22o_1 _329_ (.A1(_116_),
    .A2(_103_),
    .B1(_079_),
    .B2(_082_),
    .X(net20));
 sky130_fd_sc_hd__a21oi_1 _330_ (.A1(_111_),
    .A2(net2),
    .B1(_157_),
    .Y(_083_));
 sky130_fd_sc_hd__o22a_1 _331_ (.A1(_111_),
    .A2(net2),
    .B1(_155_),
    .B2(_083_),
    .X(_084_));
 sky130_fd_sc_hd__and2b_1 _332_ (.A_N(_118_),
    .B(_115_),
    .X(_085_));
 sky130_fd_sc_hd__nand2_1 _333_ (.A(_085_),
    .B(_117_),
    .Y(_086_));
 sky130_fd_sc_hd__o21a_1 _334_ (.A1(_085_),
    .A2(_117_),
    .B1(_129_),
    .X(_087_));
 sky130_fd_sc_hd__a21o_1 _335_ (.A1(_111_),
    .A2(net1),
    .B1(_132_),
    .X(_088_));
 sky130_fd_sc_hd__and3b_1 _336_ (.A_N(_137_),
    .B(_151_),
    .C(_088_),
    .X(_089_));
 sky130_fd_sc_hd__a31o_1 _337_ (.A1(_111_),
    .A2(net2),
    .A3(_153_),
    .B1(_089_),
    .X(_090_));
 sky130_fd_sc_hd__a211o_1 _338_ (.A1(_086_),
    .A2(_087_),
    .B1(_090_),
    .C1(_102_),
    .X(_091_));
 sky130_fd_sc_hd__o2bb2a_1 _339_ (.A1_N(net2),
    .A2_N(_103_),
    .B1(_084_),
    .B2(_091_),
    .X(net21));
 sky130_fd_sc_hd__o21ai_1 _340_ (.A1(_119_),
    .A2(_120_),
    .B1(_129_),
    .Y(_092_));
 sky130_fd_sc_hd__nor2_1 _341_ (.A(_121_),
    .B(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__or2_1 _342_ (.A(_136_),
    .B(_137_),
    .X(_094_));
 sky130_fd_sc_hd__and2b_1 _343_ (.A_N(_138_),
    .B(_151_),
    .X(_095_));
 sky130_fd_sc_hd__a21oi_1 _344_ (.A1(_105_),
    .A2(_104_),
    .B1(_157_),
    .Y(_096_));
 sky130_fd_sc_hd__o22a_1 _345_ (.A1(_105_),
    .A2(_104_),
    .B1(_155_),
    .B2(_096_),
    .X(_097_));
 sky130_fd_sc_hd__a311o_1 _346_ (.A1(_105_),
    .A2(_104_),
    .A3(_153_),
    .B1(_097_),
    .C1(_102_),
    .X(_098_));
 sky130_fd_sc_hd__a21o_1 _347_ (.A1(_094_),
    .A2(_095_),
    .B1(_098_),
    .X(_099_));
 sky130_fd_sc_hd__o2bb2a_1 _348_ (.A1_N(_104_),
    .A2_N(_103_),
    .B1(_093_),
    .B2(_099_),
    .X(net22));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_87 ();
 sky130_fd_sc_hd__buf_2 input1 (.A(A[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(A[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(A[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(A[3]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(A[4]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(A[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(A[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(A[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(B[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(B[1]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(B[2]),
    .X(net11));
 sky130_fd_sc_hd__dlymetal6s2s_1 input12 (.A(B[3]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(B[4]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(B[5]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(B[6]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(B[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(opcode[0]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(opcode[1]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(opcode[2]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(out[0]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(out[1]));
 sky130_fd_sc_hd__buf_2 output22 (.A(net22),
    .X(out[2]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(out[3]));
 sky130_fd_sc_hd__buf_2 output24 (.A(net24),
    .X(out[4]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(out[5]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(out[6]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(out[7]));
 sky130_fd_sc_hd__buf_4 output28 (.A(net28),
    .X(out[8]));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer1 (.A(_106_),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(net29),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(net29),
    .X(net31));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_113 ();
endmodule
