magic
tech sky130A
magscale 1 2
timestamp 1749470100
<< viali >>
rect 9781 17153 9815 17187
rect 10425 17153 10459 17187
rect 1409 11781 1443 11815
rect 1409 11101 1443 11135
rect 1409 10421 1443 10455
rect 18521 10421 18555 10455
rect 1409 10013 1443 10047
rect 1409 8993 1443 9027
rect 1409 8381 1443 8415
rect 9781 2397 9815 2431
rect 10425 2397 10459 2431
<< metal1 >>
rect 1104 17434 18860 17456
rect 1104 17382 2210 17434
rect 2262 17382 2274 17434
rect 2326 17382 2338 17434
rect 2390 17382 2402 17434
rect 2454 17382 2466 17434
rect 2518 17382 6210 17434
rect 6262 17382 6274 17434
rect 6326 17382 6338 17434
rect 6390 17382 6402 17434
rect 6454 17382 6466 17434
rect 6518 17382 10210 17434
rect 10262 17382 10274 17434
rect 10326 17382 10338 17434
rect 10390 17382 10402 17434
rect 10454 17382 10466 17434
rect 10518 17382 14210 17434
rect 14262 17382 14274 17434
rect 14326 17382 14338 17434
rect 14390 17382 14402 17434
rect 14454 17382 14466 17434
rect 14518 17382 18210 17434
rect 18262 17382 18274 17434
rect 18326 17382 18338 17434
rect 18390 17382 18402 17434
rect 18454 17382 18466 17434
rect 18518 17382 18860 17434
rect 1104 17360 18860 17382
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 9732 17156 9781 17184
rect 9732 17144 9738 17156
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 10134 17144 10140 17196
rect 10192 17184 10198 17196
rect 10413 17187 10471 17193
rect 10413 17184 10425 17187
rect 10192 17156 10425 17184
rect 10192 17144 10198 17156
rect 10413 17153 10425 17156
rect 10459 17153 10471 17187
rect 10413 17147 10471 17153
rect 1104 16890 18860 16912
rect 1104 16838 1550 16890
rect 1602 16838 1614 16890
rect 1666 16838 1678 16890
rect 1730 16838 1742 16890
rect 1794 16838 1806 16890
rect 1858 16838 5550 16890
rect 5602 16838 5614 16890
rect 5666 16838 5678 16890
rect 5730 16838 5742 16890
rect 5794 16838 5806 16890
rect 5858 16838 9550 16890
rect 9602 16838 9614 16890
rect 9666 16838 9678 16890
rect 9730 16838 9742 16890
rect 9794 16838 9806 16890
rect 9858 16838 13550 16890
rect 13602 16838 13614 16890
rect 13666 16838 13678 16890
rect 13730 16838 13742 16890
rect 13794 16838 13806 16890
rect 13858 16838 17550 16890
rect 17602 16838 17614 16890
rect 17666 16838 17678 16890
rect 17730 16838 17742 16890
rect 17794 16838 17806 16890
rect 17858 16838 18860 16890
rect 1104 16816 18860 16838
rect 1104 16346 18860 16368
rect 1104 16294 2210 16346
rect 2262 16294 2274 16346
rect 2326 16294 2338 16346
rect 2390 16294 2402 16346
rect 2454 16294 2466 16346
rect 2518 16294 6210 16346
rect 6262 16294 6274 16346
rect 6326 16294 6338 16346
rect 6390 16294 6402 16346
rect 6454 16294 6466 16346
rect 6518 16294 10210 16346
rect 10262 16294 10274 16346
rect 10326 16294 10338 16346
rect 10390 16294 10402 16346
rect 10454 16294 10466 16346
rect 10518 16294 14210 16346
rect 14262 16294 14274 16346
rect 14326 16294 14338 16346
rect 14390 16294 14402 16346
rect 14454 16294 14466 16346
rect 14518 16294 18210 16346
rect 18262 16294 18274 16346
rect 18326 16294 18338 16346
rect 18390 16294 18402 16346
rect 18454 16294 18466 16346
rect 18518 16294 18860 16346
rect 1104 16272 18860 16294
rect 1104 15802 18860 15824
rect 1104 15750 1550 15802
rect 1602 15750 1614 15802
rect 1666 15750 1678 15802
rect 1730 15750 1742 15802
rect 1794 15750 1806 15802
rect 1858 15750 5550 15802
rect 5602 15750 5614 15802
rect 5666 15750 5678 15802
rect 5730 15750 5742 15802
rect 5794 15750 5806 15802
rect 5858 15750 9550 15802
rect 9602 15750 9614 15802
rect 9666 15750 9678 15802
rect 9730 15750 9742 15802
rect 9794 15750 9806 15802
rect 9858 15750 13550 15802
rect 13602 15750 13614 15802
rect 13666 15750 13678 15802
rect 13730 15750 13742 15802
rect 13794 15750 13806 15802
rect 13858 15750 17550 15802
rect 17602 15750 17614 15802
rect 17666 15750 17678 15802
rect 17730 15750 17742 15802
rect 17794 15750 17806 15802
rect 17858 15750 18860 15802
rect 1104 15728 18860 15750
rect 1104 15258 18860 15280
rect 1104 15206 2210 15258
rect 2262 15206 2274 15258
rect 2326 15206 2338 15258
rect 2390 15206 2402 15258
rect 2454 15206 2466 15258
rect 2518 15206 6210 15258
rect 6262 15206 6274 15258
rect 6326 15206 6338 15258
rect 6390 15206 6402 15258
rect 6454 15206 6466 15258
rect 6518 15206 10210 15258
rect 10262 15206 10274 15258
rect 10326 15206 10338 15258
rect 10390 15206 10402 15258
rect 10454 15206 10466 15258
rect 10518 15206 14210 15258
rect 14262 15206 14274 15258
rect 14326 15206 14338 15258
rect 14390 15206 14402 15258
rect 14454 15206 14466 15258
rect 14518 15206 18210 15258
rect 18262 15206 18274 15258
rect 18326 15206 18338 15258
rect 18390 15206 18402 15258
rect 18454 15206 18466 15258
rect 18518 15206 18860 15258
rect 1104 15184 18860 15206
rect 1104 14714 18860 14736
rect 1104 14662 1550 14714
rect 1602 14662 1614 14714
rect 1666 14662 1678 14714
rect 1730 14662 1742 14714
rect 1794 14662 1806 14714
rect 1858 14662 5550 14714
rect 5602 14662 5614 14714
rect 5666 14662 5678 14714
rect 5730 14662 5742 14714
rect 5794 14662 5806 14714
rect 5858 14662 9550 14714
rect 9602 14662 9614 14714
rect 9666 14662 9678 14714
rect 9730 14662 9742 14714
rect 9794 14662 9806 14714
rect 9858 14662 13550 14714
rect 13602 14662 13614 14714
rect 13666 14662 13678 14714
rect 13730 14662 13742 14714
rect 13794 14662 13806 14714
rect 13858 14662 17550 14714
rect 17602 14662 17614 14714
rect 17666 14662 17678 14714
rect 17730 14662 17742 14714
rect 17794 14662 17806 14714
rect 17858 14662 18860 14714
rect 1104 14640 18860 14662
rect 1104 14170 18860 14192
rect 1104 14118 2210 14170
rect 2262 14118 2274 14170
rect 2326 14118 2338 14170
rect 2390 14118 2402 14170
rect 2454 14118 2466 14170
rect 2518 14118 6210 14170
rect 6262 14118 6274 14170
rect 6326 14118 6338 14170
rect 6390 14118 6402 14170
rect 6454 14118 6466 14170
rect 6518 14118 10210 14170
rect 10262 14118 10274 14170
rect 10326 14118 10338 14170
rect 10390 14118 10402 14170
rect 10454 14118 10466 14170
rect 10518 14118 14210 14170
rect 14262 14118 14274 14170
rect 14326 14118 14338 14170
rect 14390 14118 14402 14170
rect 14454 14118 14466 14170
rect 14518 14118 18210 14170
rect 18262 14118 18274 14170
rect 18326 14118 18338 14170
rect 18390 14118 18402 14170
rect 18454 14118 18466 14170
rect 18518 14118 18860 14170
rect 1104 14096 18860 14118
rect 1104 13626 18860 13648
rect 1104 13574 1550 13626
rect 1602 13574 1614 13626
rect 1666 13574 1678 13626
rect 1730 13574 1742 13626
rect 1794 13574 1806 13626
rect 1858 13574 5550 13626
rect 5602 13574 5614 13626
rect 5666 13574 5678 13626
rect 5730 13574 5742 13626
rect 5794 13574 5806 13626
rect 5858 13574 9550 13626
rect 9602 13574 9614 13626
rect 9666 13574 9678 13626
rect 9730 13574 9742 13626
rect 9794 13574 9806 13626
rect 9858 13574 13550 13626
rect 13602 13574 13614 13626
rect 13666 13574 13678 13626
rect 13730 13574 13742 13626
rect 13794 13574 13806 13626
rect 13858 13574 17550 13626
rect 17602 13574 17614 13626
rect 17666 13574 17678 13626
rect 17730 13574 17742 13626
rect 17794 13574 17806 13626
rect 17858 13574 18860 13626
rect 1104 13552 18860 13574
rect 1104 13082 18860 13104
rect 1104 13030 2210 13082
rect 2262 13030 2274 13082
rect 2326 13030 2338 13082
rect 2390 13030 2402 13082
rect 2454 13030 2466 13082
rect 2518 13030 6210 13082
rect 6262 13030 6274 13082
rect 6326 13030 6338 13082
rect 6390 13030 6402 13082
rect 6454 13030 6466 13082
rect 6518 13030 10210 13082
rect 10262 13030 10274 13082
rect 10326 13030 10338 13082
rect 10390 13030 10402 13082
rect 10454 13030 10466 13082
rect 10518 13030 14210 13082
rect 14262 13030 14274 13082
rect 14326 13030 14338 13082
rect 14390 13030 14402 13082
rect 14454 13030 14466 13082
rect 14518 13030 18210 13082
rect 18262 13030 18274 13082
rect 18326 13030 18338 13082
rect 18390 13030 18402 13082
rect 18454 13030 18466 13082
rect 18518 13030 18860 13082
rect 1104 13008 18860 13030
rect 1104 12538 18860 12560
rect 1104 12486 1550 12538
rect 1602 12486 1614 12538
rect 1666 12486 1678 12538
rect 1730 12486 1742 12538
rect 1794 12486 1806 12538
rect 1858 12486 5550 12538
rect 5602 12486 5614 12538
rect 5666 12486 5678 12538
rect 5730 12486 5742 12538
rect 5794 12486 5806 12538
rect 5858 12486 9550 12538
rect 9602 12486 9614 12538
rect 9666 12486 9678 12538
rect 9730 12486 9742 12538
rect 9794 12486 9806 12538
rect 9858 12486 13550 12538
rect 13602 12486 13614 12538
rect 13666 12486 13678 12538
rect 13730 12486 13742 12538
rect 13794 12486 13806 12538
rect 13858 12486 17550 12538
rect 17602 12486 17614 12538
rect 17666 12486 17678 12538
rect 17730 12486 17742 12538
rect 17794 12486 17806 12538
rect 17858 12486 18860 12538
rect 1104 12464 18860 12486
rect 1104 11994 18860 12016
rect 1104 11942 2210 11994
rect 2262 11942 2274 11994
rect 2326 11942 2338 11994
rect 2390 11942 2402 11994
rect 2454 11942 2466 11994
rect 2518 11942 6210 11994
rect 6262 11942 6274 11994
rect 6326 11942 6338 11994
rect 6390 11942 6402 11994
rect 6454 11942 6466 11994
rect 6518 11942 10210 11994
rect 10262 11942 10274 11994
rect 10326 11942 10338 11994
rect 10390 11942 10402 11994
rect 10454 11942 10466 11994
rect 10518 11942 14210 11994
rect 14262 11942 14274 11994
rect 14326 11942 14338 11994
rect 14390 11942 14402 11994
rect 14454 11942 14466 11994
rect 14518 11942 18210 11994
rect 18262 11942 18274 11994
rect 18326 11942 18338 11994
rect 18390 11942 18402 11994
rect 18454 11942 18466 11994
rect 18518 11942 18860 11994
rect 1104 11920 18860 11942
rect 842 11772 848 11824
rect 900 11812 906 11824
rect 1397 11815 1455 11821
rect 1397 11812 1409 11815
rect 900 11784 1409 11812
rect 900 11772 906 11784
rect 1397 11781 1409 11784
rect 1443 11781 1455 11815
rect 1397 11775 1455 11781
rect 1104 11450 18860 11472
rect 1104 11398 1550 11450
rect 1602 11398 1614 11450
rect 1666 11398 1678 11450
rect 1730 11398 1742 11450
rect 1794 11398 1806 11450
rect 1858 11398 5550 11450
rect 5602 11398 5614 11450
rect 5666 11398 5678 11450
rect 5730 11398 5742 11450
rect 5794 11398 5806 11450
rect 5858 11398 9550 11450
rect 9602 11398 9614 11450
rect 9666 11398 9678 11450
rect 9730 11398 9742 11450
rect 9794 11398 9806 11450
rect 9858 11398 13550 11450
rect 13602 11398 13614 11450
rect 13666 11398 13678 11450
rect 13730 11398 13742 11450
rect 13794 11398 13806 11450
rect 13858 11398 17550 11450
rect 17602 11398 17614 11450
rect 17666 11398 17678 11450
rect 17730 11398 17742 11450
rect 17794 11398 17806 11450
rect 17858 11398 18860 11450
rect 1104 11376 18860 11398
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 1104 10906 18860 10928
rect 1104 10854 2210 10906
rect 2262 10854 2274 10906
rect 2326 10854 2338 10906
rect 2390 10854 2402 10906
rect 2454 10854 2466 10906
rect 2518 10854 6210 10906
rect 6262 10854 6274 10906
rect 6326 10854 6338 10906
rect 6390 10854 6402 10906
rect 6454 10854 6466 10906
rect 6518 10854 10210 10906
rect 10262 10854 10274 10906
rect 10326 10854 10338 10906
rect 10390 10854 10402 10906
rect 10454 10854 10466 10906
rect 10518 10854 14210 10906
rect 14262 10854 14274 10906
rect 14326 10854 14338 10906
rect 14390 10854 14402 10906
rect 14454 10854 14466 10906
rect 14518 10854 18210 10906
rect 18262 10854 18274 10906
rect 18326 10854 18338 10906
rect 18390 10854 18402 10906
rect 18454 10854 18466 10906
rect 18518 10854 18860 10906
rect 1104 10832 18860 10854
rect 842 10412 848 10464
rect 900 10452 906 10464
rect 1397 10455 1455 10461
rect 1397 10452 1409 10455
rect 900 10424 1409 10452
rect 900 10412 906 10424
rect 1397 10421 1409 10424
rect 1443 10421 1455 10455
rect 1397 10415 1455 10421
rect 18506 10412 18512 10464
rect 18564 10412 18570 10464
rect 1104 10362 18860 10384
rect 1104 10310 1550 10362
rect 1602 10310 1614 10362
rect 1666 10310 1678 10362
rect 1730 10310 1742 10362
rect 1794 10310 1806 10362
rect 1858 10310 5550 10362
rect 5602 10310 5614 10362
rect 5666 10310 5678 10362
rect 5730 10310 5742 10362
rect 5794 10310 5806 10362
rect 5858 10310 9550 10362
rect 9602 10310 9614 10362
rect 9666 10310 9678 10362
rect 9730 10310 9742 10362
rect 9794 10310 9806 10362
rect 9858 10310 13550 10362
rect 13602 10310 13614 10362
rect 13666 10310 13678 10362
rect 13730 10310 13742 10362
rect 13794 10310 13806 10362
rect 13858 10310 17550 10362
rect 17602 10310 17614 10362
rect 17666 10310 17678 10362
rect 17730 10310 17742 10362
rect 17794 10310 17806 10362
rect 17858 10310 18860 10362
rect 1104 10288 18860 10310
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1104 9818 18860 9840
rect 1104 9766 2210 9818
rect 2262 9766 2274 9818
rect 2326 9766 2338 9818
rect 2390 9766 2402 9818
rect 2454 9766 2466 9818
rect 2518 9766 6210 9818
rect 6262 9766 6274 9818
rect 6326 9766 6338 9818
rect 6390 9766 6402 9818
rect 6454 9766 6466 9818
rect 6518 9766 10210 9818
rect 10262 9766 10274 9818
rect 10326 9766 10338 9818
rect 10390 9766 10402 9818
rect 10454 9766 10466 9818
rect 10518 9766 14210 9818
rect 14262 9766 14274 9818
rect 14326 9766 14338 9818
rect 14390 9766 14402 9818
rect 14454 9766 14466 9818
rect 14518 9766 18210 9818
rect 18262 9766 18274 9818
rect 18326 9766 18338 9818
rect 18390 9766 18402 9818
rect 18454 9766 18466 9818
rect 18518 9766 18860 9818
rect 1104 9744 18860 9766
rect 1104 9274 18860 9296
rect 1104 9222 1550 9274
rect 1602 9222 1614 9274
rect 1666 9222 1678 9274
rect 1730 9222 1742 9274
rect 1794 9222 1806 9274
rect 1858 9222 5550 9274
rect 5602 9222 5614 9274
rect 5666 9222 5678 9274
rect 5730 9222 5742 9274
rect 5794 9222 5806 9274
rect 5858 9222 9550 9274
rect 9602 9222 9614 9274
rect 9666 9222 9678 9274
rect 9730 9222 9742 9274
rect 9794 9222 9806 9274
rect 9858 9222 13550 9274
rect 13602 9222 13614 9274
rect 13666 9222 13678 9274
rect 13730 9222 13742 9274
rect 13794 9222 13806 9274
rect 13858 9222 17550 9274
rect 17602 9222 17614 9274
rect 17666 9222 17678 9274
rect 17730 9222 17742 9274
rect 17794 9222 17806 9274
rect 17858 9222 18860 9274
rect 1104 9200 18860 9222
rect 842 8984 848 9036
rect 900 9024 906 9036
rect 1397 9027 1455 9033
rect 1397 9024 1409 9027
rect 900 8996 1409 9024
rect 900 8984 906 8996
rect 1397 8993 1409 8996
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 1104 8730 18860 8752
rect 1104 8678 2210 8730
rect 2262 8678 2274 8730
rect 2326 8678 2338 8730
rect 2390 8678 2402 8730
rect 2454 8678 2466 8730
rect 2518 8678 6210 8730
rect 6262 8678 6274 8730
rect 6326 8678 6338 8730
rect 6390 8678 6402 8730
rect 6454 8678 6466 8730
rect 6518 8678 10210 8730
rect 10262 8678 10274 8730
rect 10326 8678 10338 8730
rect 10390 8678 10402 8730
rect 10454 8678 10466 8730
rect 10518 8678 14210 8730
rect 14262 8678 14274 8730
rect 14326 8678 14338 8730
rect 14390 8678 14402 8730
rect 14454 8678 14466 8730
rect 14518 8678 18210 8730
rect 18262 8678 18274 8730
rect 18326 8678 18338 8730
rect 18390 8678 18402 8730
rect 18454 8678 18466 8730
rect 18518 8678 18860 8730
rect 1104 8656 18860 8678
rect 1394 8372 1400 8424
rect 1452 8372 1458 8424
rect 1104 8186 18860 8208
rect 1104 8134 1550 8186
rect 1602 8134 1614 8186
rect 1666 8134 1678 8186
rect 1730 8134 1742 8186
rect 1794 8134 1806 8186
rect 1858 8134 5550 8186
rect 5602 8134 5614 8186
rect 5666 8134 5678 8186
rect 5730 8134 5742 8186
rect 5794 8134 5806 8186
rect 5858 8134 9550 8186
rect 9602 8134 9614 8186
rect 9666 8134 9678 8186
rect 9730 8134 9742 8186
rect 9794 8134 9806 8186
rect 9858 8134 13550 8186
rect 13602 8134 13614 8186
rect 13666 8134 13678 8186
rect 13730 8134 13742 8186
rect 13794 8134 13806 8186
rect 13858 8134 17550 8186
rect 17602 8134 17614 8186
rect 17666 8134 17678 8186
rect 17730 8134 17742 8186
rect 17794 8134 17806 8186
rect 17858 8134 18860 8186
rect 1104 8112 18860 8134
rect 1104 7642 18860 7664
rect 1104 7590 2210 7642
rect 2262 7590 2274 7642
rect 2326 7590 2338 7642
rect 2390 7590 2402 7642
rect 2454 7590 2466 7642
rect 2518 7590 6210 7642
rect 6262 7590 6274 7642
rect 6326 7590 6338 7642
rect 6390 7590 6402 7642
rect 6454 7590 6466 7642
rect 6518 7590 10210 7642
rect 10262 7590 10274 7642
rect 10326 7590 10338 7642
rect 10390 7590 10402 7642
rect 10454 7590 10466 7642
rect 10518 7590 14210 7642
rect 14262 7590 14274 7642
rect 14326 7590 14338 7642
rect 14390 7590 14402 7642
rect 14454 7590 14466 7642
rect 14518 7590 18210 7642
rect 18262 7590 18274 7642
rect 18326 7590 18338 7642
rect 18390 7590 18402 7642
rect 18454 7590 18466 7642
rect 18518 7590 18860 7642
rect 1104 7568 18860 7590
rect 1104 7098 18860 7120
rect 1104 7046 1550 7098
rect 1602 7046 1614 7098
rect 1666 7046 1678 7098
rect 1730 7046 1742 7098
rect 1794 7046 1806 7098
rect 1858 7046 5550 7098
rect 5602 7046 5614 7098
rect 5666 7046 5678 7098
rect 5730 7046 5742 7098
rect 5794 7046 5806 7098
rect 5858 7046 9550 7098
rect 9602 7046 9614 7098
rect 9666 7046 9678 7098
rect 9730 7046 9742 7098
rect 9794 7046 9806 7098
rect 9858 7046 13550 7098
rect 13602 7046 13614 7098
rect 13666 7046 13678 7098
rect 13730 7046 13742 7098
rect 13794 7046 13806 7098
rect 13858 7046 17550 7098
rect 17602 7046 17614 7098
rect 17666 7046 17678 7098
rect 17730 7046 17742 7098
rect 17794 7046 17806 7098
rect 17858 7046 18860 7098
rect 1104 7024 18860 7046
rect 1104 6554 18860 6576
rect 1104 6502 2210 6554
rect 2262 6502 2274 6554
rect 2326 6502 2338 6554
rect 2390 6502 2402 6554
rect 2454 6502 2466 6554
rect 2518 6502 6210 6554
rect 6262 6502 6274 6554
rect 6326 6502 6338 6554
rect 6390 6502 6402 6554
rect 6454 6502 6466 6554
rect 6518 6502 10210 6554
rect 10262 6502 10274 6554
rect 10326 6502 10338 6554
rect 10390 6502 10402 6554
rect 10454 6502 10466 6554
rect 10518 6502 14210 6554
rect 14262 6502 14274 6554
rect 14326 6502 14338 6554
rect 14390 6502 14402 6554
rect 14454 6502 14466 6554
rect 14518 6502 18210 6554
rect 18262 6502 18274 6554
rect 18326 6502 18338 6554
rect 18390 6502 18402 6554
rect 18454 6502 18466 6554
rect 18518 6502 18860 6554
rect 1104 6480 18860 6502
rect 1104 6010 18860 6032
rect 1104 5958 1550 6010
rect 1602 5958 1614 6010
rect 1666 5958 1678 6010
rect 1730 5958 1742 6010
rect 1794 5958 1806 6010
rect 1858 5958 5550 6010
rect 5602 5958 5614 6010
rect 5666 5958 5678 6010
rect 5730 5958 5742 6010
rect 5794 5958 5806 6010
rect 5858 5958 9550 6010
rect 9602 5958 9614 6010
rect 9666 5958 9678 6010
rect 9730 5958 9742 6010
rect 9794 5958 9806 6010
rect 9858 5958 13550 6010
rect 13602 5958 13614 6010
rect 13666 5958 13678 6010
rect 13730 5958 13742 6010
rect 13794 5958 13806 6010
rect 13858 5958 17550 6010
rect 17602 5958 17614 6010
rect 17666 5958 17678 6010
rect 17730 5958 17742 6010
rect 17794 5958 17806 6010
rect 17858 5958 18860 6010
rect 1104 5936 18860 5958
rect 1104 5466 18860 5488
rect 1104 5414 2210 5466
rect 2262 5414 2274 5466
rect 2326 5414 2338 5466
rect 2390 5414 2402 5466
rect 2454 5414 2466 5466
rect 2518 5414 6210 5466
rect 6262 5414 6274 5466
rect 6326 5414 6338 5466
rect 6390 5414 6402 5466
rect 6454 5414 6466 5466
rect 6518 5414 10210 5466
rect 10262 5414 10274 5466
rect 10326 5414 10338 5466
rect 10390 5414 10402 5466
rect 10454 5414 10466 5466
rect 10518 5414 14210 5466
rect 14262 5414 14274 5466
rect 14326 5414 14338 5466
rect 14390 5414 14402 5466
rect 14454 5414 14466 5466
rect 14518 5414 18210 5466
rect 18262 5414 18274 5466
rect 18326 5414 18338 5466
rect 18390 5414 18402 5466
rect 18454 5414 18466 5466
rect 18518 5414 18860 5466
rect 1104 5392 18860 5414
rect 1104 4922 18860 4944
rect 1104 4870 1550 4922
rect 1602 4870 1614 4922
rect 1666 4870 1678 4922
rect 1730 4870 1742 4922
rect 1794 4870 1806 4922
rect 1858 4870 5550 4922
rect 5602 4870 5614 4922
rect 5666 4870 5678 4922
rect 5730 4870 5742 4922
rect 5794 4870 5806 4922
rect 5858 4870 9550 4922
rect 9602 4870 9614 4922
rect 9666 4870 9678 4922
rect 9730 4870 9742 4922
rect 9794 4870 9806 4922
rect 9858 4870 13550 4922
rect 13602 4870 13614 4922
rect 13666 4870 13678 4922
rect 13730 4870 13742 4922
rect 13794 4870 13806 4922
rect 13858 4870 17550 4922
rect 17602 4870 17614 4922
rect 17666 4870 17678 4922
rect 17730 4870 17742 4922
rect 17794 4870 17806 4922
rect 17858 4870 18860 4922
rect 1104 4848 18860 4870
rect 1104 4378 18860 4400
rect 1104 4326 2210 4378
rect 2262 4326 2274 4378
rect 2326 4326 2338 4378
rect 2390 4326 2402 4378
rect 2454 4326 2466 4378
rect 2518 4326 6210 4378
rect 6262 4326 6274 4378
rect 6326 4326 6338 4378
rect 6390 4326 6402 4378
rect 6454 4326 6466 4378
rect 6518 4326 10210 4378
rect 10262 4326 10274 4378
rect 10326 4326 10338 4378
rect 10390 4326 10402 4378
rect 10454 4326 10466 4378
rect 10518 4326 14210 4378
rect 14262 4326 14274 4378
rect 14326 4326 14338 4378
rect 14390 4326 14402 4378
rect 14454 4326 14466 4378
rect 14518 4326 18210 4378
rect 18262 4326 18274 4378
rect 18326 4326 18338 4378
rect 18390 4326 18402 4378
rect 18454 4326 18466 4378
rect 18518 4326 18860 4378
rect 1104 4304 18860 4326
rect 1104 3834 18860 3856
rect 1104 3782 1550 3834
rect 1602 3782 1614 3834
rect 1666 3782 1678 3834
rect 1730 3782 1742 3834
rect 1794 3782 1806 3834
rect 1858 3782 5550 3834
rect 5602 3782 5614 3834
rect 5666 3782 5678 3834
rect 5730 3782 5742 3834
rect 5794 3782 5806 3834
rect 5858 3782 9550 3834
rect 9602 3782 9614 3834
rect 9666 3782 9678 3834
rect 9730 3782 9742 3834
rect 9794 3782 9806 3834
rect 9858 3782 13550 3834
rect 13602 3782 13614 3834
rect 13666 3782 13678 3834
rect 13730 3782 13742 3834
rect 13794 3782 13806 3834
rect 13858 3782 17550 3834
rect 17602 3782 17614 3834
rect 17666 3782 17678 3834
rect 17730 3782 17742 3834
rect 17794 3782 17806 3834
rect 17858 3782 18860 3834
rect 1104 3760 18860 3782
rect 1104 3290 18860 3312
rect 1104 3238 2210 3290
rect 2262 3238 2274 3290
rect 2326 3238 2338 3290
rect 2390 3238 2402 3290
rect 2454 3238 2466 3290
rect 2518 3238 6210 3290
rect 6262 3238 6274 3290
rect 6326 3238 6338 3290
rect 6390 3238 6402 3290
rect 6454 3238 6466 3290
rect 6518 3238 10210 3290
rect 10262 3238 10274 3290
rect 10326 3238 10338 3290
rect 10390 3238 10402 3290
rect 10454 3238 10466 3290
rect 10518 3238 14210 3290
rect 14262 3238 14274 3290
rect 14326 3238 14338 3290
rect 14390 3238 14402 3290
rect 14454 3238 14466 3290
rect 14518 3238 18210 3290
rect 18262 3238 18274 3290
rect 18326 3238 18338 3290
rect 18390 3238 18402 3290
rect 18454 3238 18466 3290
rect 18518 3238 18860 3290
rect 1104 3216 18860 3238
rect 1104 2746 18860 2768
rect 1104 2694 1550 2746
rect 1602 2694 1614 2746
rect 1666 2694 1678 2746
rect 1730 2694 1742 2746
rect 1794 2694 1806 2746
rect 1858 2694 5550 2746
rect 5602 2694 5614 2746
rect 5666 2694 5678 2746
rect 5730 2694 5742 2746
rect 5794 2694 5806 2746
rect 5858 2694 9550 2746
rect 9602 2694 9614 2746
rect 9666 2694 9678 2746
rect 9730 2694 9742 2746
rect 9794 2694 9806 2746
rect 9858 2694 13550 2746
rect 13602 2694 13614 2746
rect 13666 2694 13678 2746
rect 13730 2694 13742 2746
rect 13794 2694 13806 2746
rect 13858 2694 17550 2746
rect 17602 2694 17614 2746
rect 17666 2694 17678 2746
rect 17730 2694 17742 2746
rect 17794 2694 17806 2746
rect 17858 2694 18860 2746
rect 1104 2672 18860 2694
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 10134 2388 10140 2440
rect 10192 2428 10198 2440
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10192 2400 10425 2428
rect 10192 2388 10198 2400
rect 10413 2397 10425 2400
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 1104 2202 18860 2224
rect 1104 2150 2210 2202
rect 2262 2150 2274 2202
rect 2326 2150 2338 2202
rect 2390 2150 2402 2202
rect 2454 2150 2466 2202
rect 2518 2150 6210 2202
rect 6262 2150 6274 2202
rect 6326 2150 6338 2202
rect 6390 2150 6402 2202
rect 6454 2150 6466 2202
rect 6518 2150 10210 2202
rect 10262 2150 10274 2202
rect 10326 2150 10338 2202
rect 10390 2150 10402 2202
rect 10454 2150 10466 2202
rect 10518 2150 14210 2202
rect 14262 2150 14274 2202
rect 14326 2150 14338 2202
rect 14390 2150 14402 2202
rect 14454 2150 14466 2202
rect 14518 2150 18210 2202
rect 18262 2150 18274 2202
rect 18326 2150 18338 2202
rect 18390 2150 18402 2202
rect 18454 2150 18466 2202
rect 18518 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 2210 17382 2262 17434
rect 2274 17382 2326 17434
rect 2338 17382 2390 17434
rect 2402 17382 2454 17434
rect 2466 17382 2518 17434
rect 6210 17382 6262 17434
rect 6274 17382 6326 17434
rect 6338 17382 6390 17434
rect 6402 17382 6454 17434
rect 6466 17382 6518 17434
rect 10210 17382 10262 17434
rect 10274 17382 10326 17434
rect 10338 17382 10390 17434
rect 10402 17382 10454 17434
rect 10466 17382 10518 17434
rect 14210 17382 14262 17434
rect 14274 17382 14326 17434
rect 14338 17382 14390 17434
rect 14402 17382 14454 17434
rect 14466 17382 14518 17434
rect 18210 17382 18262 17434
rect 18274 17382 18326 17434
rect 18338 17382 18390 17434
rect 18402 17382 18454 17434
rect 18466 17382 18518 17434
rect 9680 17144 9732 17196
rect 10140 17144 10192 17196
rect 1550 16838 1602 16890
rect 1614 16838 1666 16890
rect 1678 16838 1730 16890
rect 1742 16838 1794 16890
rect 1806 16838 1858 16890
rect 5550 16838 5602 16890
rect 5614 16838 5666 16890
rect 5678 16838 5730 16890
rect 5742 16838 5794 16890
rect 5806 16838 5858 16890
rect 9550 16838 9602 16890
rect 9614 16838 9666 16890
rect 9678 16838 9730 16890
rect 9742 16838 9794 16890
rect 9806 16838 9858 16890
rect 13550 16838 13602 16890
rect 13614 16838 13666 16890
rect 13678 16838 13730 16890
rect 13742 16838 13794 16890
rect 13806 16838 13858 16890
rect 17550 16838 17602 16890
rect 17614 16838 17666 16890
rect 17678 16838 17730 16890
rect 17742 16838 17794 16890
rect 17806 16838 17858 16890
rect 2210 16294 2262 16346
rect 2274 16294 2326 16346
rect 2338 16294 2390 16346
rect 2402 16294 2454 16346
rect 2466 16294 2518 16346
rect 6210 16294 6262 16346
rect 6274 16294 6326 16346
rect 6338 16294 6390 16346
rect 6402 16294 6454 16346
rect 6466 16294 6518 16346
rect 10210 16294 10262 16346
rect 10274 16294 10326 16346
rect 10338 16294 10390 16346
rect 10402 16294 10454 16346
rect 10466 16294 10518 16346
rect 14210 16294 14262 16346
rect 14274 16294 14326 16346
rect 14338 16294 14390 16346
rect 14402 16294 14454 16346
rect 14466 16294 14518 16346
rect 18210 16294 18262 16346
rect 18274 16294 18326 16346
rect 18338 16294 18390 16346
rect 18402 16294 18454 16346
rect 18466 16294 18518 16346
rect 1550 15750 1602 15802
rect 1614 15750 1666 15802
rect 1678 15750 1730 15802
rect 1742 15750 1794 15802
rect 1806 15750 1858 15802
rect 5550 15750 5602 15802
rect 5614 15750 5666 15802
rect 5678 15750 5730 15802
rect 5742 15750 5794 15802
rect 5806 15750 5858 15802
rect 9550 15750 9602 15802
rect 9614 15750 9666 15802
rect 9678 15750 9730 15802
rect 9742 15750 9794 15802
rect 9806 15750 9858 15802
rect 13550 15750 13602 15802
rect 13614 15750 13666 15802
rect 13678 15750 13730 15802
rect 13742 15750 13794 15802
rect 13806 15750 13858 15802
rect 17550 15750 17602 15802
rect 17614 15750 17666 15802
rect 17678 15750 17730 15802
rect 17742 15750 17794 15802
rect 17806 15750 17858 15802
rect 2210 15206 2262 15258
rect 2274 15206 2326 15258
rect 2338 15206 2390 15258
rect 2402 15206 2454 15258
rect 2466 15206 2518 15258
rect 6210 15206 6262 15258
rect 6274 15206 6326 15258
rect 6338 15206 6390 15258
rect 6402 15206 6454 15258
rect 6466 15206 6518 15258
rect 10210 15206 10262 15258
rect 10274 15206 10326 15258
rect 10338 15206 10390 15258
rect 10402 15206 10454 15258
rect 10466 15206 10518 15258
rect 14210 15206 14262 15258
rect 14274 15206 14326 15258
rect 14338 15206 14390 15258
rect 14402 15206 14454 15258
rect 14466 15206 14518 15258
rect 18210 15206 18262 15258
rect 18274 15206 18326 15258
rect 18338 15206 18390 15258
rect 18402 15206 18454 15258
rect 18466 15206 18518 15258
rect 1550 14662 1602 14714
rect 1614 14662 1666 14714
rect 1678 14662 1730 14714
rect 1742 14662 1794 14714
rect 1806 14662 1858 14714
rect 5550 14662 5602 14714
rect 5614 14662 5666 14714
rect 5678 14662 5730 14714
rect 5742 14662 5794 14714
rect 5806 14662 5858 14714
rect 9550 14662 9602 14714
rect 9614 14662 9666 14714
rect 9678 14662 9730 14714
rect 9742 14662 9794 14714
rect 9806 14662 9858 14714
rect 13550 14662 13602 14714
rect 13614 14662 13666 14714
rect 13678 14662 13730 14714
rect 13742 14662 13794 14714
rect 13806 14662 13858 14714
rect 17550 14662 17602 14714
rect 17614 14662 17666 14714
rect 17678 14662 17730 14714
rect 17742 14662 17794 14714
rect 17806 14662 17858 14714
rect 2210 14118 2262 14170
rect 2274 14118 2326 14170
rect 2338 14118 2390 14170
rect 2402 14118 2454 14170
rect 2466 14118 2518 14170
rect 6210 14118 6262 14170
rect 6274 14118 6326 14170
rect 6338 14118 6390 14170
rect 6402 14118 6454 14170
rect 6466 14118 6518 14170
rect 10210 14118 10262 14170
rect 10274 14118 10326 14170
rect 10338 14118 10390 14170
rect 10402 14118 10454 14170
rect 10466 14118 10518 14170
rect 14210 14118 14262 14170
rect 14274 14118 14326 14170
rect 14338 14118 14390 14170
rect 14402 14118 14454 14170
rect 14466 14118 14518 14170
rect 18210 14118 18262 14170
rect 18274 14118 18326 14170
rect 18338 14118 18390 14170
rect 18402 14118 18454 14170
rect 18466 14118 18518 14170
rect 1550 13574 1602 13626
rect 1614 13574 1666 13626
rect 1678 13574 1730 13626
rect 1742 13574 1794 13626
rect 1806 13574 1858 13626
rect 5550 13574 5602 13626
rect 5614 13574 5666 13626
rect 5678 13574 5730 13626
rect 5742 13574 5794 13626
rect 5806 13574 5858 13626
rect 9550 13574 9602 13626
rect 9614 13574 9666 13626
rect 9678 13574 9730 13626
rect 9742 13574 9794 13626
rect 9806 13574 9858 13626
rect 13550 13574 13602 13626
rect 13614 13574 13666 13626
rect 13678 13574 13730 13626
rect 13742 13574 13794 13626
rect 13806 13574 13858 13626
rect 17550 13574 17602 13626
rect 17614 13574 17666 13626
rect 17678 13574 17730 13626
rect 17742 13574 17794 13626
rect 17806 13574 17858 13626
rect 2210 13030 2262 13082
rect 2274 13030 2326 13082
rect 2338 13030 2390 13082
rect 2402 13030 2454 13082
rect 2466 13030 2518 13082
rect 6210 13030 6262 13082
rect 6274 13030 6326 13082
rect 6338 13030 6390 13082
rect 6402 13030 6454 13082
rect 6466 13030 6518 13082
rect 10210 13030 10262 13082
rect 10274 13030 10326 13082
rect 10338 13030 10390 13082
rect 10402 13030 10454 13082
rect 10466 13030 10518 13082
rect 14210 13030 14262 13082
rect 14274 13030 14326 13082
rect 14338 13030 14390 13082
rect 14402 13030 14454 13082
rect 14466 13030 14518 13082
rect 18210 13030 18262 13082
rect 18274 13030 18326 13082
rect 18338 13030 18390 13082
rect 18402 13030 18454 13082
rect 18466 13030 18518 13082
rect 1550 12486 1602 12538
rect 1614 12486 1666 12538
rect 1678 12486 1730 12538
rect 1742 12486 1794 12538
rect 1806 12486 1858 12538
rect 5550 12486 5602 12538
rect 5614 12486 5666 12538
rect 5678 12486 5730 12538
rect 5742 12486 5794 12538
rect 5806 12486 5858 12538
rect 9550 12486 9602 12538
rect 9614 12486 9666 12538
rect 9678 12486 9730 12538
rect 9742 12486 9794 12538
rect 9806 12486 9858 12538
rect 13550 12486 13602 12538
rect 13614 12486 13666 12538
rect 13678 12486 13730 12538
rect 13742 12486 13794 12538
rect 13806 12486 13858 12538
rect 17550 12486 17602 12538
rect 17614 12486 17666 12538
rect 17678 12486 17730 12538
rect 17742 12486 17794 12538
rect 17806 12486 17858 12538
rect 2210 11942 2262 11994
rect 2274 11942 2326 11994
rect 2338 11942 2390 11994
rect 2402 11942 2454 11994
rect 2466 11942 2518 11994
rect 6210 11942 6262 11994
rect 6274 11942 6326 11994
rect 6338 11942 6390 11994
rect 6402 11942 6454 11994
rect 6466 11942 6518 11994
rect 10210 11942 10262 11994
rect 10274 11942 10326 11994
rect 10338 11942 10390 11994
rect 10402 11942 10454 11994
rect 10466 11942 10518 11994
rect 14210 11942 14262 11994
rect 14274 11942 14326 11994
rect 14338 11942 14390 11994
rect 14402 11942 14454 11994
rect 14466 11942 14518 11994
rect 18210 11942 18262 11994
rect 18274 11942 18326 11994
rect 18338 11942 18390 11994
rect 18402 11942 18454 11994
rect 18466 11942 18518 11994
rect 848 11772 900 11824
rect 1550 11398 1602 11450
rect 1614 11398 1666 11450
rect 1678 11398 1730 11450
rect 1742 11398 1794 11450
rect 1806 11398 1858 11450
rect 5550 11398 5602 11450
rect 5614 11398 5666 11450
rect 5678 11398 5730 11450
rect 5742 11398 5794 11450
rect 5806 11398 5858 11450
rect 9550 11398 9602 11450
rect 9614 11398 9666 11450
rect 9678 11398 9730 11450
rect 9742 11398 9794 11450
rect 9806 11398 9858 11450
rect 13550 11398 13602 11450
rect 13614 11398 13666 11450
rect 13678 11398 13730 11450
rect 13742 11398 13794 11450
rect 13806 11398 13858 11450
rect 17550 11398 17602 11450
rect 17614 11398 17666 11450
rect 17678 11398 17730 11450
rect 17742 11398 17794 11450
rect 17806 11398 17858 11450
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2210 10854 2262 10906
rect 2274 10854 2326 10906
rect 2338 10854 2390 10906
rect 2402 10854 2454 10906
rect 2466 10854 2518 10906
rect 6210 10854 6262 10906
rect 6274 10854 6326 10906
rect 6338 10854 6390 10906
rect 6402 10854 6454 10906
rect 6466 10854 6518 10906
rect 10210 10854 10262 10906
rect 10274 10854 10326 10906
rect 10338 10854 10390 10906
rect 10402 10854 10454 10906
rect 10466 10854 10518 10906
rect 14210 10854 14262 10906
rect 14274 10854 14326 10906
rect 14338 10854 14390 10906
rect 14402 10854 14454 10906
rect 14466 10854 14518 10906
rect 18210 10854 18262 10906
rect 18274 10854 18326 10906
rect 18338 10854 18390 10906
rect 18402 10854 18454 10906
rect 18466 10854 18518 10906
rect 848 10412 900 10464
rect 18512 10455 18564 10464
rect 18512 10421 18521 10455
rect 18521 10421 18555 10455
rect 18555 10421 18564 10455
rect 18512 10412 18564 10421
rect 1550 10310 1602 10362
rect 1614 10310 1666 10362
rect 1678 10310 1730 10362
rect 1742 10310 1794 10362
rect 1806 10310 1858 10362
rect 5550 10310 5602 10362
rect 5614 10310 5666 10362
rect 5678 10310 5730 10362
rect 5742 10310 5794 10362
rect 5806 10310 5858 10362
rect 9550 10310 9602 10362
rect 9614 10310 9666 10362
rect 9678 10310 9730 10362
rect 9742 10310 9794 10362
rect 9806 10310 9858 10362
rect 13550 10310 13602 10362
rect 13614 10310 13666 10362
rect 13678 10310 13730 10362
rect 13742 10310 13794 10362
rect 13806 10310 13858 10362
rect 17550 10310 17602 10362
rect 17614 10310 17666 10362
rect 17678 10310 17730 10362
rect 17742 10310 17794 10362
rect 17806 10310 17858 10362
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2210 9766 2262 9818
rect 2274 9766 2326 9818
rect 2338 9766 2390 9818
rect 2402 9766 2454 9818
rect 2466 9766 2518 9818
rect 6210 9766 6262 9818
rect 6274 9766 6326 9818
rect 6338 9766 6390 9818
rect 6402 9766 6454 9818
rect 6466 9766 6518 9818
rect 10210 9766 10262 9818
rect 10274 9766 10326 9818
rect 10338 9766 10390 9818
rect 10402 9766 10454 9818
rect 10466 9766 10518 9818
rect 14210 9766 14262 9818
rect 14274 9766 14326 9818
rect 14338 9766 14390 9818
rect 14402 9766 14454 9818
rect 14466 9766 14518 9818
rect 18210 9766 18262 9818
rect 18274 9766 18326 9818
rect 18338 9766 18390 9818
rect 18402 9766 18454 9818
rect 18466 9766 18518 9818
rect 1550 9222 1602 9274
rect 1614 9222 1666 9274
rect 1678 9222 1730 9274
rect 1742 9222 1794 9274
rect 1806 9222 1858 9274
rect 5550 9222 5602 9274
rect 5614 9222 5666 9274
rect 5678 9222 5730 9274
rect 5742 9222 5794 9274
rect 5806 9222 5858 9274
rect 9550 9222 9602 9274
rect 9614 9222 9666 9274
rect 9678 9222 9730 9274
rect 9742 9222 9794 9274
rect 9806 9222 9858 9274
rect 13550 9222 13602 9274
rect 13614 9222 13666 9274
rect 13678 9222 13730 9274
rect 13742 9222 13794 9274
rect 13806 9222 13858 9274
rect 17550 9222 17602 9274
rect 17614 9222 17666 9274
rect 17678 9222 17730 9274
rect 17742 9222 17794 9274
rect 17806 9222 17858 9274
rect 848 8984 900 9036
rect 2210 8678 2262 8730
rect 2274 8678 2326 8730
rect 2338 8678 2390 8730
rect 2402 8678 2454 8730
rect 2466 8678 2518 8730
rect 6210 8678 6262 8730
rect 6274 8678 6326 8730
rect 6338 8678 6390 8730
rect 6402 8678 6454 8730
rect 6466 8678 6518 8730
rect 10210 8678 10262 8730
rect 10274 8678 10326 8730
rect 10338 8678 10390 8730
rect 10402 8678 10454 8730
rect 10466 8678 10518 8730
rect 14210 8678 14262 8730
rect 14274 8678 14326 8730
rect 14338 8678 14390 8730
rect 14402 8678 14454 8730
rect 14466 8678 14518 8730
rect 18210 8678 18262 8730
rect 18274 8678 18326 8730
rect 18338 8678 18390 8730
rect 18402 8678 18454 8730
rect 18466 8678 18518 8730
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 1550 8134 1602 8186
rect 1614 8134 1666 8186
rect 1678 8134 1730 8186
rect 1742 8134 1794 8186
rect 1806 8134 1858 8186
rect 5550 8134 5602 8186
rect 5614 8134 5666 8186
rect 5678 8134 5730 8186
rect 5742 8134 5794 8186
rect 5806 8134 5858 8186
rect 9550 8134 9602 8186
rect 9614 8134 9666 8186
rect 9678 8134 9730 8186
rect 9742 8134 9794 8186
rect 9806 8134 9858 8186
rect 13550 8134 13602 8186
rect 13614 8134 13666 8186
rect 13678 8134 13730 8186
rect 13742 8134 13794 8186
rect 13806 8134 13858 8186
rect 17550 8134 17602 8186
rect 17614 8134 17666 8186
rect 17678 8134 17730 8186
rect 17742 8134 17794 8186
rect 17806 8134 17858 8186
rect 2210 7590 2262 7642
rect 2274 7590 2326 7642
rect 2338 7590 2390 7642
rect 2402 7590 2454 7642
rect 2466 7590 2518 7642
rect 6210 7590 6262 7642
rect 6274 7590 6326 7642
rect 6338 7590 6390 7642
rect 6402 7590 6454 7642
rect 6466 7590 6518 7642
rect 10210 7590 10262 7642
rect 10274 7590 10326 7642
rect 10338 7590 10390 7642
rect 10402 7590 10454 7642
rect 10466 7590 10518 7642
rect 14210 7590 14262 7642
rect 14274 7590 14326 7642
rect 14338 7590 14390 7642
rect 14402 7590 14454 7642
rect 14466 7590 14518 7642
rect 18210 7590 18262 7642
rect 18274 7590 18326 7642
rect 18338 7590 18390 7642
rect 18402 7590 18454 7642
rect 18466 7590 18518 7642
rect 1550 7046 1602 7098
rect 1614 7046 1666 7098
rect 1678 7046 1730 7098
rect 1742 7046 1794 7098
rect 1806 7046 1858 7098
rect 5550 7046 5602 7098
rect 5614 7046 5666 7098
rect 5678 7046 5730 7098
rect 5742 7046 5794 7098
rect 5806 7046 5858 7098
rect 9550 7046 9602 7098
rect 9614 7046 9666 7098
rect 9678 7046 9730 7098
rect 9742 7046 9794 7098
rect 9806 7046 9858 7098
rect 13550 7046 13602 7098
rect 13614 7046 13666 7098
rect 13678 7046 13730 7098
rect 13742 7046 13794 7098
rect 13806 7046 13858 7098
rect 17550 7046 17602 7098
rect 17614 7046 17666 7098
rect 17678 7046 17730 7098
rect 17742 7046 17794 7098
rect 17806 7046 17858 7098
rect 2210 6502 2262 6554
rect 2274 6502 2326 6554
rect 2338 6502 2390 6554
rect 2402 6502 2454 6554
rect 2466 6502 2518 6554
rect 6210 6502 6262 6554
rect 6274 6502 6326 6554
rect 6338 6502 6390 6554
rect 6402 6502 6454 6554
rect 6466 6502 6518 6554
rect 10210 6502 10262 6554
rect 10274 6502 10326 6554
rect 10338 6502 10390 6554
rect 10402 6502 10454 6554
rect 10466 6502 10518 6554
rect 14210 6502 14262 6554
rect 14274 6502 14326 6554
rect 14338 6502 14390 6554
rect 14402 6502 14454 6554
rect 14466 6502 14518 6554
rect 18210 6502 18262 6554
rect 18274 6502 18326 6554
rect 18338 6502 18390 6554
rect 18402 6502 18454 6554
rect 18466 6502 18518 6554
rect 1550 5958 1602 6010
rect 1614 5958 1666 6010
rect 1678 5958 1730 6010
rect 1742 5958 1794 6010
rect 1806 5958 1858 6010
rect 5550 5958 5602 6010
rect 5614 5958 5666 6010
rect 5678 5958 5730 6010
rect 5742 5958 5794 6010
rect 5806 5958 5858 6010
rect 9550 5958 9602 6010
rect 9614 5958 9666 6010
rect 9678 5958 9730 6010
rect 9742 5958 9794 6010
rect 9806 5958 9858 6010
rect 13550 5958 13602 6010
rect 13614 5958 13666 6010
rect 13678 5958 13730 6010
rect 13742 5958 13794 6010
rect 13806 5958 13858 6010
rect 17550 5958 17602 6010
rect 17614 5958 17666 6010
rect 17678 5958 17730 6010
rect 17742 5958 17794 6010
rect 17806 5958 17858 6010
rect 2210 5414 2262 5466
rect 2274 5414 2326 5466
rect 2338 5414 2390 5466
rect 2402 5414 2454 5466
rect 2466 5414 2518 5466
rect 6210 5414 6262 5466
rect 6274 5414 6326 5466
rect 6338 5414 6390 5466
rect 6402 5414 6454 5466
rect 6466 5414 6518 5466
rect 10210 5414 10262 5466
rect 10274 5414 10326 5466
rect 10338 5414 10390 5466
rect 10402 5414 10454 5466
rect 10466 5414 10518 5466
rect 14210 5414 14262 5466
rect 14274 5414 14326 5466
rect 14338 5414 14390 5466
rect 14402 5414 14454 5466
rect 14466 5414 14518 5466
rect 18210 5414 18262 5466
rect 18274 5414 18326 5466
rect 18338 5414 18390 5466
rect 18402 5414 18454 5466
rect 18466 5414 18518 5466
rect 1550 4870 1602 4922
rect 1614 4870 1666 4922
rect 1678 4870 1730 4922
rect 1742 4870 1794 4922
rect 1806 4870 1858 4922
rect 5550 4870 5602 4922
rect 5614 4870 5666 4922
rect 5678 4870 5730 4922
rect 5742 4870 5794 4922
rect 5806 4870 5858 4922
rect 9550 4870 9602 4922
rect 9614 4870 9666 4922
rect 9678 4870 9730 4922
rect 9742 4870 9794 4922
rect 9806 4870 9858 4922
rect 13550 4870 13602 4922
rect 13614 4870 13666 4922
rect 13678 4870 13730 4922
rect 13742 4870 13794 4922
rect 13806 4870 13858 4922
rect 17550 4870 17602 4922
rect 17614 4870 17666 4922
rect 17678 4870 17730 4922
rect 17742 4870 17794 4922
rect 17806 4870 17858 4922
rect 2210 4326 2262 4378
rect 2274 4326 2326 4378
rect 2338 4326 2390 4378
rect 2402 4326 2454 4378
rect 2466 4326 2518 4378
rect 6210 4326 6262 4378
rect 6274 4326 6326 4378
rect 6338 4326 6390 4378
rect 6402 4326 6454 4378
rect 6466 4326 6518 4378
rect 10210 4326 10262 4378
rect 10274 4326 10326 4378
rect 10338 4326 10390 4378
rect 10402 4326 10454 4378
rect 10466 4326 10518 4378
rect 14210 4326 14262 4378
rect 14274 4326 14326 4378
rect 14338 4326 14390 4378
rect 14402 4326 14454 4378
rect 14466 4326 14518 4378
rect 18210 4326 18262 4378
rect 18274 4326 18326 4378
rect 18338 4326 18390 4378
rect 18402 4326 18454 4378
rect 18466 4326 18518 4378
rect 1550 3782 1602 3834
rect 1614 3782 1666 3834
rect 1678 3782 1730 3834
rect 1742 3782 1794 3834
rect 1806 3782 1858 3834
rect 5550 3782 5602 3834
rect 5614 3782 5666 3834
rect 5678 3782 5730 3834
rect 5742 3782 5794 3834
rect 5806 3782 5858 3834
rect 9550 3782 9602 3834
rect 9614 3782 9666 3834
rect 9678 3782 9730 3834
rect 9742 3782 9794 3834
rect 9806 3782 9858 3834
rect 13550 3782 13602 3834
rect 13614 3782 13666 3834
rect 13678 3782 13730 3834
rect 13742 3782 13794 3834
rect 13806 3782 13858 3834
rect 17550 3782 17602 3834
rect 17614 3782 17666 3834
rect 17678 3782 17730 3834
rect 17742 3782 17794 3834
rect 17806 3782 17858 3834
rect 2210 3238 2262 3290
rect 2274 3238 2326 3290
rect 2338 3238 2390 3290
rect 2402 3238 2454 3290
rect 2466 3238 2518 3290
rect 6210 3238 6262 3290
rect 6274 3238 6326 3290
rect 6338 3238 6390 3290
rect 6402 3238 6454 3290
rect 6466 3238 6518 3290
rect 10210 3238 10262 3290
rect 10274 3238 10326 3290
rect 10338 3238 10390 3290
rect 10402 3238 10454 3290
rect 10466 3238 10518 3290
rect 14210 3238 14262 3290
rect 14274 3238 14326 3290
rect 14338 3238 14390 3290
rect 14402 3238 14454 3290
rect 14466 3238 14518 3290
rect 18210 3238 18262 3290
rect 18274 3238 18326 3290
rect 18338 3238 18390 3290
rect 18402 3238 18454 3290
rect 18466 3238 18518 3290
rect 1550 2694 1602 2746
rect 1614 2694 1666 2746
rect 1678 2694 1730 2746
rect 1742 2694 1794 2746
rect 1806 2694 1858 2746
rect 5550 2694 5602 2746
rect 5614 2694 5666 2746
rect 5678 2694 5730 2746
rect 5742 2694 5794 2746
rect 5806 2694 5858 2746
rect 9550 2694 9602 2746
rect 9614 2694 9666 2746
rect 9678 2694 9730 2746
rect 9742 2694 9794 2746
rect 9806 2694 9858 2746
rect 13550 2694 13602 2746
rect 13614 2694 13666 2746
rect 13678 2694 13730 2746
rect 13742 2694 13794 2746
rect 13806 2694 13858 2746
rect 17550 2694 17602 2746
rect 17614 2694 17666 2746
rect 17678 2694 17730 2746
rect 17742 2694 17794 2746
rect 17806 2694 17858 2746
rect 9680 2388 9732 2440
rect 10140 2388 10192 2440
rect 2210 2150 2262 2202
rect 2274 2150 2326 2202
rect 2338 2150 2390 2202
rect 2402 2150 2454 2202
rect 2466 2150 2518 2202
rect 6210 2150 6262 2202
rect 6274 2150 6326 2202
rect 6338 2150 6390 2202
rect 6402 2150 6454 2202
rect 6466 2150 6518 2202
rect 10210 2150 10262 2202
rect 10274 2150 10326 2202
rect 10338 2150 10390 2202
rect 10402 2150 10454 2202
rect 10466 2150 10518 2202
rect 14210 2150 14262 2202
rect 14274 2150 14326 2202
rect 14338 2150 14390 2202
rect 14402 2150 14454 2202
rect 14466 2150 14518 2202
rect 18210 2150 18262 2202
rect 18274 2150 18326 2202
rect 18338 2150 18390 2202
rect 18402 2150 18454 2202
rect 18466 2150 18518 2202
<< metal2 >>
rect 9678 19200 9734 20000
rect 10322 19200 10378 20000
rect 2210 17436 2518 17445
rect 2210 17434 2216 17436
rect 2272 17434 2296 17436
rect 2352 17434 2376 17436
rect 2432 17434 2456 17436
rect 2512 17434 2518 17436
rect 2272 17382 2274 17434
rect 2454 17382 2456 17434
rect 2210 17380 2216 17382
rect 2272 17380 2296 17382
rect 2352 17380 2376 17382
rect 2432 17380 2456 17382
rect 2512 17380 2518 17382
rect 2210 17371 2518 17380
rect 6210 17436 6518 17445
rect 6210 17434 6216 17436
rect 6272 17434 6296 17436
rect 6352 17434 6376 17436
rect 6432 17434 6456 17436
rect 6512 17434 6518 17436
rect 6272 17382 6274 17434
rect 6454 17382 6456 17434
rect 6210 17380 6216 17382
rect 6272 17380 6296 17382
rect 6352 17380 6376 17382
rect 6432 17380 6456 17382
rect 6512 17380 6518 17382
rect 6210 17371 6518 17380
rect 9692 17202 9720 19200
rect 10336 17626 10364 19200
rect 10152 17598 10364 17626
rect 10152 17202 10180 17598
rect 10210 17436 10518 17445
rect 10210 17434 10216 17436
rect 10272 17434 10296 17436
rect 10352 17434 10376 17436
rect 10432 17434 10456 17436
rect 10512 17434 10518 17436
rect 10272 17382 10274 17434
rect 10454 17382 10456 17434
rect 10210 17380 10216 17382
rect 10272 17380 10296 17382
rect 10352 17380 10376 17382
rect 10432 17380 10456 17382
rect 10512 17380 10518 17382
rect 10210 17371 10518 17380
rect 14210 17436 14518 17445
rect 14210 17434 14216 17436
rect 14272 17434 14296 17436
rect 14352 17434 14376 17436
rect 14432 17434 14456 17436
rect 14512 17434 14518 17436
rect 14272 17382 14274 17434
rect 14454 17382 14456 17434
rect 14210 17380 14216 17382
rect 14272 17380 14296 17382
rect 14352 17380 14376 17382
rect 14432 17380 14456 17382
rect 14512 17380 14518 17382
rect 14210 17371 14518 17380
rect 18210 17436 18518 17445
rect 18210 17434 18216 17436
rect 18272 17434 18296 17436
rect 18352 17434 18376 17436
rect 18432 17434 18456 17436
rect 18512 17434 18518 17436
rect 18272 17382 18274 17434
rect 18454 17382 18456 17434
rect 18210 17380 18216 17382
rect 18272 17380 18296 17382
rect 18352 17380 18376 17382
rect 18432 17380 18456 17382
rect 18512 17380 18518 17382
rect 18210 17371 18518 17380
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 1550 16892 1858 16901
rect 1550 16890 1556 16892
rect 1612 16890 1636 16892
rect 1692 16890 1716 16892
rect 1772 16890 1796 16892
rect 1852 16890 1858 16892
rect 1612 16838 1614 16890
rect 1794 16838 1796 16890
rect 1550 16836 1556 16838
rect 1612 16836 1636 16838
rect 1692 16836 1716 16838
rect 1772 16836 1796 16838
rect 1852 16836 1858 16838
rect 1550 16827 1858 16836
rect 5550 16892 5858 16901
rect 5550 16890 5556 16892
rect 5612 16890 5636 16892
rect 5692 16890 5716 16892
rect 5772 16890 5796 16892
rect 5852 16890 5858 16892
rect 5612 16838 5614 16890
rect 5794 16838 5796 16890
rect 5550 16836 5556 16838
rect 5612 16836 5636 16838
rect 5692 16836 5716 16838
rect 5772 16836 5796 16838
rect 5852 16836 5858 16838
rect 5550 16827 5858 16836
rect 9550 16892 9858 16901
rect 9550 16890 9556 16892
rect 9612 16890 9636 16892
rect 9692 16890 9716 16892
rect 9772 16890 9796 16892
rect 9852 16890 9858 16892
rect 9612 16838 9614 16890
rect 9794 16838 9796 16890
rect 9550 16836 9556 16838
rect 9612 16836 9636 16838
rect 9692 16836 9716 16838
rect 9772 16836 9796 16838
rect 9852 16836 9858 16838
rect 9550 16827 9858 16836
rect 13550 16892 13858 16901
rect 13550 16890 13556 16892
rect 13612 16890 13636 16892
rect 13692 16890 13716 16892
rect 13772 16890 13796 16892
rect 13852 16890 13858 16892
rect 13612 16838 13614 16890
rect 13794 16838 13796 16890
rect 13550 16836 13556 16838
rect 13612 16836 13636 16838
rect 13692 16836 13716 16838
rect 13772 16836 13796 16838
rect 13852 16836 13858 16838
rect 13550 16827 13858 16836
rect 17550 16892 17858 16901
rect 17550 16890 17556 16892
rect 17612 16890 17636 16892
rect 17692 16890 17716 16892
rect 17772 16890 17796 16892
rect 17852 16890 17858 16892
rect 17612 16838 17614 16890
rect 17794 16838 17796 16890
rect 17550 16836 17556 16838
rect 17612 16836 17636 16838
rect 17692 16836 17716 16838
rect 17772 16836 17796 16838
rect 17852 16836 17858 16838
rect 17550 16827 17858 16836
rect 2210 16348 2518 16357
rect 2210 16346 2216 16348
rect 2272 16346 2296 16348
rect 2352 16346 2376 16348
rect 2432 16346 2456 16348
rect 2512 16346 2518 16348
rect 2272 16294 2274 16346
rect 2454 16294 2456 16346
rect 2210 16292 2216 16294
rect 2272 16292 2296 16294
rect 2352 16292 2376 16294
rect 2432 16292 2456 16294
rect 2512 16292 2518 16294
rect 2210 16283 2518 16292
rect 6210 16348 6518 16357
rect 6210 16346 6216 16348
rect 6272 16346 6296 16348
rect 6352 16346 6376 16348
rect 6432 16346 6456 16348
rect 6512 16346 6518 16348
rect 6272 16294 6274 16346
rect 6454 16294 6456 16346
rect 6210 16292 6216 16294
rect 6272 16292 6296 16294
rect 6352 16292 6376 16294
rect 6432 16292 6456 16294
rect 6512 16292 6518 16294
rect 6210 16283 6518 16292
rect 10210 16348 10518 16357
rect 10210 16346 10216 16348
rect 10272 16346 10296 16348
rect 10352 16346 10376 16348
rect 10432 16346 10456 16348
rect 10512 16346 10518 16348
rect 10272 16294 10274 16346
rect 10454 16294 10456 16346
rect 10210 16292 10216 16294
rect 10272 16292 10296 16294
rect 10352 16292 10376 16294
rect 10432 16292 10456 16294
rect 10512 16292 10518 16294
rect 10210 16283 10518 16292
rect 14210 16348 14518 16357
rect 14210 16346 14216 16348
rect 14272 16346 14296 16348
rect 14352 16346 14376 16348
rect 14432 16346 14456 16348
rect 14512 16346 14518 16348
rect 14272 16294 14274 16346
rect 14454 16294 14456 16346
rect 14210 16292 14216 16294
rect 14272 16292 14296 16294
rect 14352 16292 14376 16294
rect 14432 16292 14456 16294
rect 14512 16292 14518 16294
rect 14210 16283 14518 16292
rect 18210 16348 18518 16357
rect 18210 16346 18216 16348
rect 18272 16346 18296 16348
rect 18352 16346 18376 16348
rect 18432 16346 18456 16348
rect 18512 16346 18518 16348
rect 18272 16294 18274 16346
rect 18454 16294 18456 16346
rect 18210 16292 18216 16294
rect 18272 16292 18296 16294
rect 18352 16292 18376 16294
rect 18432 16292 18456 16294
rect 18512 16292 18518 16294
rect 18210 16283 18518 16292
rect 1550 15804 1858 15813
rect 1550 15802 1556 15804
rect 1612 15802 1636 15804
rect 1692 15802 1716 15804
rect 1772 15802 1796 15804
rect 1852 15802 1858 15804
rect 1612 15750 1614 15802
rect 1794 15750 1796 15802
rect 1550 15748 1556 15750
rect 1612 15748 1636 15750
rect 1692 15748 1716 15750
rect 1772 15748 1796 15750
rect 1852 15748 1858 15750
rect 1550 15739 1858 15748
rect 5550 15804 5858 15813
rect 5550 15802 5556 15804
rect 5612 15802 5636 15804
rect 5692 15802 5716 15804
rect 5772 15802 5796 15804
rect 5852 15802 5858 15804
rect 5612 15750 5614 15802
rect 5794 15750 5796 15802
rect 5550 15748 5556 15750
rect 5612 15748 5636 15750
rect 5692 15748 5716 15750
rect 5772 15748 5796 15750
rect 5852 15748 5858 15750
rect 5550 15739 5858 15748
rect 9550 15804 9858 15813
rect 9550 15802 9556 15804
rect 9612 15802 9636 15804
rect 9692 15802 9716 15804
rect 9772 15802 9796 15804
rect 9852 15802 9858 15804
rect 9612 15750 9614 15802
rect 9794 15750 9796 15802
rect 9550 15748 9556 15750
rect 9612 15748 9636 15750
rect 9692 15748 9716 15750
rect 9772 15748 9796 15750
rect 9852 15748 9858 15750
rect 9550 15739 9858 15748
rect 13550 15804 13858 15813
rect 13550 15802 13556 15804
rect 13612 15802 13636 15804
rect 13692 15802 13716 15804
rect 13772 15802 13796 15804
rect 13852 15802 13858 15804
rect 13612 15750 13614 15802
rect 13794 15750 13796 15802
rect 13550 15748 13556 15750
rect 13612 15748 13636 15750
rect 13692 15748 13716 15750
rect 13772 15748 13796 15750
rect 13852 15748 13858 15750
rect 13550 15739 13858 15748
rect 17550 15804 17858 15813
rect 17550 15802 17556 15804
rect 17612 15802 17636 15804
rect 17692 15802 17716 15804
rect 17772 15802 17796 15804
rect 17852 15802 17858 15804
rect 17612 15750 17614 15802
rect 17794 15750 17796 15802
rect 17550 15748 17556 15750
rect 17612 15748 17636 15750
rect 17692 15748 17716 15750
rect 17772 15748 17796 15750
rect 17852 15748 17858 15750
rect 17550 15739 17858 15748
rect 2210 15260 2518 15269
rect 2210 15258 2216 15260
rect 2272 15258 2296 15260
rect 2352 15258 2376 15260
rect 2432 15258 2456 15260
rect 2512 15258 2518 15260
rect 2272 15206 2274 15258
rect 2454 15206 2456 15258
rect 2210 15204 2216 15206
rect 2272 15204 2296 15206
rect 2352 15204 2376 15206
rect 2432 15204 2456 15206
rect 2512 15204 2518 15206
rect 2210 15195 2518 15204
rect 6210 15260 6518 15269
rect 6210 15258 6216 15260
rect 6272 15258 6296 15260
rect 6352 15258 6376 15260
rect 6432 15258 6456 15260
rect 6512 15258 6518 15260
rect 6272 15206 6274 15258
rect 6454 15206 6456 15258
rect 6210 15204 6216 15206
rect 6272 15204 6296 15206
rect 6352 15204 6376 15206
rect 6432 15204 6456 15206
rect 6512 15204 6518 15206
rect 6210 15195 6518 15204
rect 10210 15260 10518 15269
rect 10210 15258 10216 15260
rect 10272 15258 10296 15260
rect 10352 15258 10376 15260
rect 10432 15258 10456 15260
rect 10512 15258 10518 15260
rect 10272 15206 10274 15258
rect 10454 15206 10456 15258
rect 10210 15204 10216 15206
rect 10272 15204 10296 15206
rect 10352 15204 10376 15206
rect 10432 15204 10456 15206
rect 10512 15204 10518 15206
rect 10210 15195 10518 15204
rect 14210 15260 14518 15269
rect 14210 15258 14216 15260
rect 14272 15258 14296 15260
rect 14352 15258 14376 15260
rect 14432 15258 14456 15260
rect 14512 15258 14518 15260
rect 14272 15206 14274 15258
rect 14454 15206 14456 15258
rect 14210 15204 14216 15206
rect 14272 15204 14296 15206
rect 14352 15204 14376 15206
rect 14432 15204 14456 15206
rect 14512 15204 14518 15206
rect 14210 15195 14518 15204
rect 18210 15260 18518 15269
rect 18210 15258 18216 15260
rect 18272 15258 18296 15260
rect 18352 15258 18376 15260
rect 18432 15258 18456 15260
rect 18512 15258 18518 15260
rect 18272 15206 18274 15258
rect 18454 15206 18456 15258
rect 18210 15204 18216 15206
rect 18272 15204 18296 15206
rect 18352 15204 18376 15206
rect 18432 15204 18456 15206
rect 18512 15204 18518 15206
rect 18210 15195 18518 15204
rect 1550 14716 1858 14725
rect 1550 14714 1556 14716
rect 1612 14714 1636 14716
rect 1692 14714 1716 14716
rect 1772 14714 1796 14716
rect 1852 14714 1858 14716
rect 1612 14662 1614 14714
rect 1794 14662 1796 14714
rect 1550 14660 1556 14662
rect 1612 14660 1636 14662
rect 1692 14660 1716 14662
rect 1772 14660 1796 14662
rect 1852 14660 1858 14662
rect 1550 14651 1858 14660
rect 5550 14716 5858 14725
rect 5550 14714 5556 14716
rect 5612 14714 5636 14716
rect 5692 14714 5716 14716
rect 5772 14714 5796 14716
rect 5852 14714 5858 14716
rect 5612 14662 5614 14714
rect 5794 14662 5796 14714
rect 5550 14660 5556 14662
rect 5612 14660 5636 14662
rect 5692 14660 5716 14662
rect 5772 14660 5796 14662
rect 5852 14660 5858 14662
rect 5550 14651 5858 14660
rect 9550 14716 9858 14725
rect 9550 14714 9556 14716
rect 9612 14714 9636 14716
rect 9692 14714 9716 14716
rect 9772 14714 9796 14716
rect 9852 14714 9858 14716
rect 9612 14662 9614 14714
rect 9794 14662 9796 14714
rect 9550 14660 9556 14662
rect 9612 14660 9636 14662
rect 9692 14660 9716 14662
rect 9772 14660 9796 14662
rect 9852 14660 9858 14662
rect 9550 14651 9858 14660
rect 13550 14716 13858 14725
rect 13550 14714 13556 14716
rect 13612 14714 13636 14716
rect 13692 14714 13716 14716
rect 13772 14714 13796 14716
rect 13852 14714 13858 14716
rect 13612 14662 13614 14714
rect 13794 14662 13796 14714
rect 13550 14660 13556 14662
rect 13612 14660 13636 14662
rect 13692 14660 13716 14662
rect 13772 14660 13796 14662
rect 13852 14660 13858 14662
rect 13550 14651 13858 14660
rect 17550 14716 17858 14725
rect 17550 14714 17556 14716
rect 17612 14714 17636 14716
rect 17692 14714 17716 14716
rect 17772 14714 17796 14716
rect 17852 14714 17858 14716
rect 17612 14662 17614 14714
rect 17794 14662 17796 14714
rect 17550 14660 17556 14662
rect 17612 14660 17636 14662
rect 17692 14660 17716 14662
rect 17772 14660 17796 14662
rect 17852 14660 17858 14662
rect 17550 14651 17858 14660
rect 2210 14172 2518 14181
rect 2210 14170 2216 14172
rect 2272 14170 2296 14172
rect 2352 14170 2376 14172
rect 2432 14170 2456 14172
rect 2512 14170 2518 14172
rect 2272 14118 2274 14170
rect 2454 14118 2456 14170
rect 2210 14116 2216 14118
rect 2272 14116 2296 14118
rect 2352 14116 2376 14118
rect 2432 14116 2456 14118
rect 2512 14116 2518 14118
rect 2210 14107 2518 14116
rect 6210 14172 6518 14181
rect 6210 14170 6216 14172
rect 6272 14170 6296 14172
rect 6352 14170 6376 14172
rect 6432 14170 6456 14172
rect 6512 14170 6518 14172
rect 6272 14118 6274 14170
rect 6454 14118 6456 14170
rect 6210 14116 6216 14118
rect 6272 14116 6296 14118
rect 6352 14116 6376 14118
rect 6432 14116 6456 14118
rect 6512 14116 6518 14118
rect 6210 14107 6518 14116
rect 10210 14172 10518 14181
rect 10210 14170 10216 14172
rect 10272 14170 10296 14172
rect 10352 14170 10376 14172
rect 10432 14170 10456 14172
rect 10512 14170 10518 14172
rect 10272 14118 10274 14170
rect 10454 14118 10456 14170
rect 10210 14116 10216 14118
rect 10272 14116 10296 14118
rect 10352 14116 10376 14118
rect 10432 14116 10456 14118
rect 10512 14116 10518 14118
rect 10210 14107 10518 14116
rect 14210 14172 14518 14181
rect 14210 14170 14216 14172
rect 14272 14170 14296 14172
rect 14352 14170 14376 14172
rect 14432 14170 14456 14172
rect 14512 14170 14518 14172
rect 14272 14118 14274 14170
rect 14454 14118 14456 14170
rect 14210 14116 14216 14118
rect 14272 14116 14296 14118
rect 14352 14116 14376 14118
rect 14432 14116 14456 14118
rect 14512 14116 14518 14118
rect 14210 14107 14518 14116
rect 18210 14172 18518 14181
rect 18210 14170 18216 14172
rect 18272 14170 18296 14172
rect 18352 14170 18376 14172
rect 18432 14170 18456 14172
rect 18512 14170 18518 14172
rect 18272 14118 18274 14170
rect 18454 14118 18456 14170
rect 18210 14116 18216 14118
rect 18272 14116 18296 14118
rect 18352 14116 18376 14118
rect 18432 14116 18456 14118
rect 18512 14116 18518 14118
rect 18210 14107 18518 14116
rect 1550 13628 1858 13637
rect 1550 13626 1556 13628
rect 1612 13626 1636 13628
rect 1692 13626 1716 13628
rect 1772 13626 1796 13628
rect 1852 13626 1858 13628
rect 1612 13574 1614 13626
rect 1794 13574 1796 13626
rect 1550 13572 1556 13574
rect 1612 13572 1636 13574
rect 1692 13572 1716 13574
rect 1772 13572 1796 13574
rect 1852 13572 1858 13574
rect 1550 13563 1858 13572
rect 5550 13628 5858 13637
rect 5550 13626 5556 13628
rect 5612 13626 5636 13628
rect 5692 13626 5716 13628
rect 5772 13626 5796 13628
rect 5852 13626 5858 13628
rect 5612 13574 5614 13626
rect 5794 13574 5796 13626
rect 5550 13572 5556 13574
rect 5612 13572 5636 13574
rect 5692 13572 5716 13574
rect 5772 13572 5796 13574
rect 5852 13572 5858 13574
rect 5550 13563 5858 13572
rect 9550 13628 9858 13637
rect 9550 13626 9556 13628
rect 9612 13626 9636 13628
rect 9692 13626 9716 13628
rect 9772 13626 9796 13628
rect 9852 13626 9858 13628
rect 9612 13574 9614 13626
rect 9794 13574 9796 13626
rect 9550 13572 9556 13574
rect 9612 13572 9636 13574
rect 9692 13572 9716 13574
rect 9772 13572 9796 13574
rect 9852 13572 9858 13574
rect 9550 13563 9858 13572
rect 13550 13628 13858 13637
rect 13550 13626 13556 13628
rect 13612 13626 13636 13628
rect 13692 13626 13716 13628
rect 13772 13626 13796 13628
rect 13852 13626 13858 13628
rect 13612 13574 13614 13626
rect 13794 13574 13796 13626
rect 13550 13572 13556 13574
rect 13612 13572 13636 13574
rect 13692 13572 13716 13574
rect 13772 13572 13796 13574
rect 13852 13572 13858 13574
rect 13550 13563 13858 13572
rect 17550 13628 17858 13637
rect 17550 13626 17556 13628
rect 17612 13626 17636 13628
rect 17692 13626 17716 13628
rect 17772 13626 17796 13628
rect 17852 13626 17858 13628
rect 17612 13574 17614 13626
rect 17794 13574 17796 13626
rect 17550 13572 17556 13574
rect 17612 13572 17636 13574
rect 17692 13572 17716 13574
rect 17772 13572 17796 13574
rect 17852 13572 17858 13574
rect 17550 13563 17858 13572
rect 2210 13084 2518 13093
rect 2210 13082 2216 13084
rect 2272 13082 2296 13084
rect 2352 13082 2376 13084
rect 2432 13082 2456 13084
rect 2512 13082 2518 13084
rect 2272 13030 2274 13082
rect 2454 13030 2456 13082
rect 2210 13028 2216 13030
rect 2272 13028 2296 13030
rect 2352 13028 2376 13030
rect 2432 13028 2456 13030
rect 2512 13028 2518 13030
rect 2210 13019 2518 13028
rect 6210 13084 6518 13093
rect 6210 13082 6216 13084
rect 6272 13082 6296 13084
rect 6352 13082 6376 13084
rect 6432 13082 6456 13084
rect 6512 13082 6518 13084
rect 6272 13030 6274 13082
rect 6454 13030 6456 13082
rect 6210 13028 6216 13030
rect 6272 13028 6296 13030
rect 6352 13028 6376 13030
rect 6432 13028 6456 13030
rect 6512 13028 6518 13030
rect 6210 13019 6518 13028
rect 10210 13084 10518 13093
rect 10210 13082 10216 13084
rect 10272 13082 10296 13084
rect 10352 13082 10376 13084
rect 10432 13082 10456 13084
rect 10512 13082 10518 13084
rect 10272 13030 10274 13082
rect 10454 13030 10456 13082
rect 10210 13028 10216 13030
rect 10272 13028 10296 13030
rect 10352 13028 10376 13030
rect 10432 13028 10456 13030
rect 10512 13028 10518 13030
rect 10210 13019 10518 13028
rect 14210 13084 14518 13093
rect 14210 13082 14216 13084
rect 14272 13082 14296 13084
rect 14352 13082 14376 13084
rect 14432 13082 14456 13084
rect 14512 13082 14518 13084
rect 14272 13030 14274 13082
rect 14454 13030 14456 13082
rect 14210 13028 14216 13030
rect 14272 13028 14296 13030
rect 14352 13028 14376 13030
rect 14432 13028 14456 13030
rect 14512 13028 14518 13030
rect 14210 13019 14518 13028
rect 18210 13084 18518 13093
rect 18210 13082 18216 13084
rect 18272 13082 18296 13084
rect 18352 13082 18376 13084
rect 18432 13082 18456 13084
rect 18512 13082 18518 13084
rect 18272 13030 18274 13082
rect 18454 13030 18456 13082
rect 18210 13028 18216 13030
rect 18272 13028 18296 13030
rect 18352 13028 18376 13030
rect 18432 13028 18456 13030
rect 18512 13028 18518 13030
rect 18210 13019 18518 13028
rect 1550 12540 1858 12549
rect 1550 12538 1556 12540
rect 1612 12538 1636 12540
rect 1692 12538 1716 12540
rect 1772 12538 1796 12540
rect 1852 12538 1858 12540
rect 1612 12486 1614 12538
rect 1794 12486 1796 12538
rect 1550 12484 1556 12486
rect 1612 12484 1636 12486
rect 1692 12484 1716 12486
rect 1772 12484 1796 12486
rect 1852 12484 1858 12486
rect 1550 12475 1858 12484
rect 5550 12540 5858 12549
rect 5550 12538 5556 12540
rect 5612 12538 5636 12540
rect 5692 12538 5716 12540
rect 5772 12538 5796 12540
rect 5852 12538 5858 12540
rect 5612 12486 5614 12538
rect 5794 12486 5796 12538
rect 5550 12484 5556 12486
rect 5612 12484 5636 12486
rect 5692 12484 5716 12486
rect 5772 12484 5796 12486
rect 5852 12484 5858 12486
rect 5550 12475 5858 12484
rect 9550 12540 9858 12549
rect 9550 12538 9556 12540
rect 9612 12538 9636 12540
rect 9692 12538 9716 12540
rect 9772 12538 9796 12540
rect 9852 12538 9858 12540
rect 9612 12486 9614 12538
rect 9794 12486 9796 12538
rect 9550 12484 9556 12486
rect 9612 12484 9636 12486
rect 9692 12484 9716 12486
rect 9772 12484 9796 12486
rect 9852 12484 9858 12486
rect 9550 12475 9858 12484
rect 13550 12540 13858 12549
rect 13550 12538 13556 12540
rect 13612 12538 13636 12540
rect 13692 12538 13716 12540
rect 13772 12538 13796 12540
rect 13852 12538 13858 12540
rect 13612 12486 13614 12538
rect 13794 12486 13796 12538
rect 13550 12484 13556 12486
rect 13612 12484 13636 12486
rect 13692 12484 13716 12486
rect 13772 12484 13796 12486
rect 13852 12484 13858 12486
rect 13550 12475 13858 12484
rect 17550 12540 17858 12549
rect 17550 12538 17556 12540
rect 17612 12538 17636 12540
rect 17692 12538 17716 12540
rect 17772 12538 17796 12540
rect 17852 12538 17858 12540
rect 17612 12486 17614 12538
rect 17794 12486 17796 12538
rect 17550 12484 17556 12486
rect 17612 12484 17636 12486
rect 17692 12484 17716 12486
rect 17772 12484 17796 12486
rect 17852 12484 17858 12486
rect 17550 12475 17858 12484
rect 2210 11996 2518 12005
rect 2210 11994 2216 11996
rect 2272 11994 2296 11996
rect 2352 11994 2376 11996
rect 2432 11994 2456 11996
rect 2512 11994 2518 11996
rect 2272 11942 2274 11994
rect 2454 11942 2456 11994
rect 2210 11940 2216 11942
rect 2272 11940 2296 11942
rect 2352 11940 2376 11942
rect 2432 11940 2456 11942
rect 2512 11940 2518 11942
rect 2210 11931 2518 11940
rect 6210 11996 6518 12005
rect 6210 11994 6216 11996
rect 6272 11994 6296 11996
rect 6352 11994 6376 11996
rect 6432 11994 6456 11996
rect 6512 11994 6518 11996
rect 6272 11942 6274 11994
rect 6454 11942 6456 11994
rect 6210 11940 6216 11942
rect 6272 11940 6296 11942
rect 6352 11940 6376 11942
rect 6432 11940 6456 11942
rect 6512 11940 6518 11942
rect 6210 11931 6518 11940
rect 10210 11996 10518 12005
rect 10210 11994 10216 11996
rect 10272 11994 10296 11996
rect 10352 11994 10376 11996
rect 10432 11994 10456 11996
rect 10512 11994 10518 11996
rect 10272 11942 10274 11994
rect 10454 11942 10456 11994
rect 10210 11940 10216 11942
rect 10272 11940 10296 11942
rect 10352 11940 10376 11942
rect 10432 11940 10456 11942
rect 10512 11940 10518 11942
rect 10210 11931 10518 11940
rect 14210 11996 14518 12005
rect 14210 11994 14216 11996
rect 14272 11994 14296 11996
rect 14352 11994 14376 11996
rect 14432 11994 14456 11996
rect 14512 11994 14518 11996
rect 14272 11942 14274 11994
rect 14454 11942 14456 11994
rect 14210 11940 14216 11942
rect 14272 11940 14296 11942
rect 14352 11940 14376 11942
rect 14432 11940 14456 11942
rect 14512 11940 14518 11942
rect 14210 11931 14518 11940
rect 18210 11996 18518 12005
rect 18210 11994 18216 11996
rect 18272 11994 18296 11996
rect 18352 11994 18376 11996
rect 18432 11994 18456 11996
rect 18512 11994 18518 11996
rect 18272 11942 18274 11994
rect 18454 11942 18456 11994
rect 18210 11940 18216 11942
rect 18272 11940 18296 11942
rect 18352 11940 18376 11942
rect 18432 11940 18456 11942
rect 18512 11940 18518 11942
rect 18210 11931 18518 11940
rect 848 11824 900 11830
rect 846 11792 848 11801
rect 900 11792 902 11801
rect 846 11727 902 11736
rect 1550 11452 1858 11461
rect 1550 11450 1556 11452
rect 1612 11450 1636 11452
rect 1692 11450 1716 11452
rect 1772 11450 1796 11452
rect 1852 11450 1858 11452
rect 1612 11398 1614 11450
rect 1794 11398 1796 11450
rect 1550 11396 1556 11398
rect 1612 11396 1636 11398
rect 1692 11396 1716 11398
rect 1772 11396 1796 11398
rect 1852 11396 1858 11398
rect 1550 11387 1858 11396
rect 5550 11452 5858 11461
rect 5550 11450 5556 11452
rect 5612 11450 5636 11452
rect 5692 11450 5716 11452
rect 5772 11450 5796 11452
rect 5852 11450 5858 11452
rect 5612 11398 5614 11450
rect 5794 11398 5796 11450
rect 5550 11396 5556 11398
rect 5612 11396 5636 11398
rect 5692 11396 5716 11398
rect 5772 11396 5796 11398
rect 5852 11396 5858 11398
rect 5550 11387 5858 11396
rect 9550 11452 9858 11461
rect 9550 11450 9556 11452
rect 9612 11450 9636 11452
rect 9692 11450 9716 11452
rect 9772 11450 9796 11452
rect 9852 11450 9858 11452
rect 9612 11398 9614 11450
rect 9794 11398 9796 11450
rect 9550 11396 9556 11398
rect 9612 11396 9636 11398
rect 9692 11396 9716 11398
rect 9772 11396 9796 11398
rect 9852 11396 9858 11398
rect 9550 11387 9858 11396
rect 13550 11452 13858 11461
rect 13550 11450 13556 11452
rect 13612 11450 13636 11452
rect 13692 11450 13716 11452
rect 13772 11450 13796 11452
rect 13852 11450 13858 11452
rect 13612 11398 13614 11450
rect 13794 11398 13796 11450
rect 13550 11396 13556 11398
rect 13612 11396 13636 11398
rect 13692 11396 13716 11398
rect 13772 11396 13796 11398
rect 13852 11396 13858 11398
rect 13550 11387 13858 11396
rect 17550 11452 17858 11461
rect 17550 11450 17556 11452
rect 17612 11450 17636 11452
rect 17692 11450 17716 11452
rect 17772 11450 17796 11452
rect 17852 11450 17858 11452
rect 17612 11398 17614 11450
rect 17794 11398 17796 11450
rect 17550 11396 17556 11398
rect 17612 11396 17636 11398
rect 17692 11396 17716 11398
rect 17772 11396 17796 11398
rect 17852 11396 17858 11398
rect 17550 11387 17858 11396
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 2210 10908 2518 10917
rect 2210 10906 2216 10908
rect 2272 10906 2296 10908
rect 2352 10906 2376 10908
rect 2432 10906 2456 10908
rect 2512 10906 2518 10908
rect 2272 10854 2274 10906
rect 2454 10854 2456 10906
rect 2210 10852 2216 10854
rect 2272 10852 2296 10854
rect 2352 10852 2376 10854
rect 2432 10852 2456 10854
rect 2512 10852 2518 10854
rect 2210 10843 2518 10852
rect 6210 10908 6518 10917
rect 6210 10906 6216 10908
rect 6272 10906 6296 10908
rect 6352 10906 6376 10908
rect 6432 10906 6456 10908
rect 6512 10906 6518 10908
rect 6272 10854 6274 10906
rect 6454 10854 6456 10906
rect 6210 10852 6216 10854
rect 6272 10852 6296 10854
rect 6352 10852 6376 10854
rect 6432 10852 6456 10854
rect 6512 10852 6518 10854
rect 6210 10843 6518 10852
rect 10210 10908 10518 10917
rect 10210 10906 10216 10908
rect 10272 10906 10296 10908
rect 10352 10906 10376 10908
rect 10432 10906 10456 10908
rect 10512 10906 10518 10908
rect 10272 10854 10274 10906
rect 10454 10854 10456 10906
rect 10210 10852 10216 10854
rect 10272 10852 10296 10854
rect 10352 10852 10376 10854
rect 10432 10852 10456 10854
rect 10512 10852 10518 10854
rect 10210 10843 10518 10852
rect 14210 10908 14518 10917
rect 14210 10906 14216 10908
rect 14272 10906 14296 10908
rect 14352 10906 14376 10908
rect 14432 10906 14456 10908
rect 14512 10906 14518 10908
rect 14272 10854 14274 10906
rect 14454 10854 14456 10906
rect 14210 10852 14216 10854
rect 14272 10852 14296 10854
rect 14352 10852 14376 10854
rect 14432 10852 14456 10854
rect 14512 10852 14518 10854
rect 14210 10843 14518 10852
rect 18210 10908 18518 10917
rect 18210 10906 18216 10908
rect 18272 10906 18296 10908
rect 18352 10906 18376 10908
rect 18432 10906 18456 10908
rect 18512 10906 18518 10908
rect 18272 10854 18274 10906
rect 18454 10854 18456 10906
rect 18210 10852 18216 10854
rect 18272 10852 18296 10854
rect 18352 10852 18376 10854
rect 18432 10852 18456 10854
rect 18512 10852 18518 10854
rect 18210 10843 18518 10852
rect 848 10464 900 10470
rect 846 10432 848 10441
rect 18512 10464 18564 10470
rect 900 10432 902 10441
rect 18512 10406 18564 10412
rect 846 10367 902 10376
rect 1550 10364 1858 10373
rect 1550 10362 1556 10364
rect 1612 10362 1636 10364
rect 1692 10362 1716 10364
rect 1772 10362 1796 10364
rect 1852 10362 1858 10364
rect 1612 10310 1614 10362
rect 1794 10310 1796 10362
rect 1550 10308 1556 10310
rect 1612 10308 1636 10310
rect 1692 10308 1716 10310
rect 1772 10308 1796 10310
rect 1852 10308 1858 10310
rect 1550 10299 1858 10308
rect 5550 10364 5858 10373
rect 5550 10362 5556 10364
rect 5612 10362 5636 10364
rect 5692 10362 5716 10364
rect 5772 10362 5796 10364
rect 5852 10362 5858 10364
rect 5612 10310 5614 10362
rect 5794 10310 5796 10362
rect 5550 10308 5556 10310
rect 5612 10308 5636 10310
rect 5692 10308 5716 10310
rect 5772 10308 5796 10310
rect 5852 10308 5858 10310
rect 5550 10299 5858 10308
rect 9550 10364 9858 10373
rect 9550 10362 9556 10364
rect 9612 10362 9636 10364
rect 9692 10362 9716 10364
rect 9772 10362 9796 10364
rect 9852 10362 9858 10364
rect 9612 10310 9614 10362
rect 9794 10310 9796 10362
rect 9550 10308 9556 10310
rect 9612 10308 9636 10310
rect 9692 10308 9716 10310
rect 9772 10308 9796 10310
rect 9852 10308 9858 10310
rect 9550 10299 9858 10308
rect 13550 10364 13858 10373
rect 13550 10362 13556 10364
rect 13612 10362 13636 10364
rect 13692 10362 13716 10364
rect 13772 10362 13796 10364
rect 13852 10362 13858 10364
rect 13612 10310 13614 10362
rect 13794 10310 13796 10362
rect 13550 10308 13556 10310
rect 13612 10308 13636 10310
rect 13692 10308 13716 10310
rect 13772 10308 13796 10310
rect 13852 10308 13858 10310
rect 13550 10299 13858 10308
rect 17550 10364 17858 10373
rect 17550 10362 17556 10364
rect 17612 10362 17636 10364
rect 17692 10362 17716 10364
rect 17772 10362 17796 10364
rect 17852 10362 17858 10364
rect 17612 10310 17614 10362
rect 17794 10310 17796 10362
rect 17550 10308 17556 10310
rect 17612 10308 17636 10310
rect 17692 10308 17716 10310
rect 17772 10308 17796 10310
rect 17852 10308 17858 10310
rect 17550 10299 17858 10308
rect 18524 10305 18552 10406
rect 18510 10296 18566 10305
rect 18510 10231 18566 10240
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 2210 9820 2518 9829
rect 2210 9818 2216 9820
rect 2272 9818 2296 9820
rect 2352 9818 2376 9820
rect 2432 9818 2456 9820
rect 2512 9818 2518 9820
rect 2272 9766 2274 9818
rect 2454 9766 2456 9818
rect 2210 9764 2216 9766
rect 2272 9764 2296 9766
rect 2352 9764 2376 9766
rect 2432 9764 2456 9766
rect 2512 9764 2518 9766
rect 2210 9755 2518 9764
rect 6210 9820 6518 9829
rect 6210 9818 6216 9820
rect 6272 9818 6296 9820
rect 6352 9818 6376 9820
rect 6432 9818 6456 9820
rect 6512 9818 6518 9820
rect 6272 9766 6274 9818
rect 6454 9766 6456 9818
rect 6210 9764 6216 9766
rect 6272 9764 6296 9766
rect 6352 9764 6376 9766
rect 6432 9764 6456 9766
rect 6512 9764 6518 9766
rect 6210 9755 6518 9764
rect 10210 9820 10518 9829
rect 10210 9818 10216 9820
rect 10272 9818 10296 9820
rect 10352 9818 10376 9820
rect 10432 9818 10456 9820
rect 10512 9818 10518 9820
rect 10272 9766 10274 9818
rect 10454 9766 10456 9818
rect 10210 9764 10216 9766
rect 10272 9764 10296 9766
rect 10352 9764 10376 9766
rect 10432 9764 10456 9766
rect 10512 9764 10518 9766
rect 10210 9755 10518 9764
rect 14210 9820 14518 9829
rect 14210 9818 14216 9820
rect 14272 9818 14296 9820
rect 14352 9818 14376 9820
rect 14432 9818 14456 9820
rect 14512 9818 14518 9820
rect 14272 9766 14274 9818
rect 14454 9766 14456 9818
rect 14210 9764 14216 9766
rect 14272 9764 14296 9766
rect 14352 9764 14376 9766
rect 14432 9764 14456 9766
rect 14512 9764 14518 9766
rect 14210 9755 14518 9764
rect 18210 9820 18518 9829
rect 18210 9818 18216 9820
rect 18272 9818 18296 9820
rect 18352 9818 18376 9820
rect 18432 9818 18456 9820
rect 18512 9818 18518 9820
rect 18272 9766 18274 9818
rect 18454 9766 18456 9818
rect 18210 9764 18216 9766
rect 18272 9764 18296 9766
rect 18352 9764 18376 9766
rect 18432 9764 18456 9766
rect 18512 9764 18518 9766
rect 18210 9755 18518 9764
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1550 9276 1858 9285
rect 1550 9274 1556 9276
rect 1612 9274 1636 9276
rect 1692 9274 1716 9276
rect 1772 9274 1796 9276
rect 1852 9274 1858 9276
rect 1612 9222 1614 9274
rect 1794 9222 1796 9274
rect 1550 9220 1556 9222
rect 1612 9220 1636 9222
rect 1692 9220 1716 9222
rect 1772 9220 1796 9222
rect 1852 9220 1858 9222
rect 1550 9211 1858 9220
rect 5550 9276 5858 9285
rect 5550 9274 5556 9276
rect 5612 9274 5636 9276
rect 5692 9274 5716 9276
rect 5772 9274 5796 9276
rect 5852 9274 5858 9276
rect 5612 9222 5614 9274
rect 5794 9222 5796 9274
rect 5550 9220 5556 9222
rect 5612 9220 5636 9222
rect 5692 9220 5716 9222
rect 5772 9220 5796 9222
rect 5852 9220 5858 9222
rect 5550 9211 5858 9220
rect 9550 9276 9858 9285
rect 9550 9274 9556 9276
rect 9612 9274 9636 9276
rect 9692 9274 9716 9276
rect 9772 9274 9796 9276
rect 9852 9274 9858 9276
rect 9612 9222 9614 9274
rect 9794 9222 9796 9274
rect 9550 9220 9556 9222
rect 9612 9220 9636 9222
rect 9692 9220 9716 9222
rect 9772 9220 9796 9222
rect 9852 9220 9858 9222
rect 9550 9211 9858 9220
rect 13550 9276 13858 9285
rect 13550 9274 13556 9276
rect 13612 9274 13636 9276
rect 13692 9274 13716 9276
rect 13772 9274 13796 9276
rect 13852 9274 13858 9276
rect 13612 9222 13614 9274
rect 13794 9222 13796 9274
rect 13550 9220 13556 9222
rect 13612 9220 13636 9222
rect 13692 9220 13716 9222
rect 13772 9220 13796 9222
rect 13852 9220 13858 9222
rect 13550 9211 13858 9220
rect 17550 9276 17858 9285
rect 17550 9274 17556 9276
rect 17612 9274 17636 9276
rect 17692 9274 17716 9276
rect 17772 9274 17796 9276
rect 17852 9274 17858 9276
rect 17612 9222 17614 9274
rect 17794 9222 17796 9274
rect 17550 9220 17556 9222
rect 17612 9220 17636 9222
rect 17692 9220 17716 9222
rect 17772 9220 17796 9222
rect 17852 9220 17858 9222
rect 17550 9211 17858 9220
rect 846 9072 902 9081
rect 846 9007 848 9016
rect 900 9007 902 9016
rect 848 8978 900 8984
rect 2210 8732 2518 8741
rect 2210 8730 2216 8732
rect 2272 8730 2296 8732
rect 2352 8730 2376 8732
rect 2432 8730 2456 8732
rect 2512 8730 2518 8732
rect 2272 8678 2274 8730
rect 2454 8678 2456 8730
rect 2210 8676 2216 8678
rect 2272 8676 2296 8678
rect 2352 8676 2376 8678
rect 2432 8676 2456 8678
rect 2512 8676 2518 8678
rect 2210 8667 2518 8676
rect 6210 8732 6518 8741
rect 6210 8730 6216 8732
rect 6272 8730 6296 8732
rect 6352 8730 6376 8732
rect 6432 8730 6456 8732
rect 6512 8730 6518 8732
rect 6272 8678 6274 8730
rect 6454 8678 6456 8730
rect 6210 8676 6216 8678
rect 6272 8676 6296 8678
rect 6352 8676 6376 8678
rect 6432 8676 6456 8678
rect 6512 8676 6518 8678
rect 6210 8667 6518 8676
rect 10210 8732 10518 8741
rect 10210 8730 10216 8732
rect 10272 8730 10296 8732
rect 10352 8730 10376 8732
rect 10432 8730 10456 8732
rect 10512 8730 10518 8732
rect 10272 8678 10274 8730
rect 10454 8678 10456 8730
rect 10210 8676 10216 8678
rect 10272 8676 10296 8678
rect 10352 8676 10376 8678
rect 10432 8676 10456 8678
rect 10512 8676 10518 8678
rect 10210 8667 10518 8676
rect 14210 8732 14518 8741
rect 14210 8730 14216 8732
rect 14272 8730 14296 8732
rect 14352 8730 14376 8732
rect 14432 8730 14456 8732
rect 14512 8730 14518 8732
rect 14272 8678 14274 8730
rect 14454 8678 14456 8730
rect 14210 8676 14216 8678
rect 14272 8676 14296 8678
rect 14352 8676 14376 8678
rect 14432 8676 14456 8678
rect 14512 8676 14518 8678
rect 14210 8667 14518 8676
rect 18210 8732 18518 8741
rect 18210 8730 18216 8732
rect 18272 8730 18296 8732
rect 18352 8730 18376 8732
rect 18432 8730 18456 8732
rect 18512 8730 18518 8732
rect 18272 8678 18274 8730
rect 18454 8678 18456 8730
rect 18210 8676 18216 8678
rect 18272 8676 18296 8678
rect 18352 8676 18376 8678
rect 18432 8676 18456 8678
rect 18512 8676 18518 8678
rect 18210 8667 18518 8676
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 1550 8188 1858 8197
rect 1550 8186 1556 8188
rect 1612 8186 1636 8188
rect 1692 8186 1716 8188
rect 1772 8186 1796 8188
rect 1852 8186 1858 8188
rect 1612 8134 1614 8186
rect 1794 8134 1796 8186
rect 1550 8132 1556 8134
rect 1612 8132 1636 8134
rect 1692 8132 1716 8134
rect 1772 8132 1796 8134
rect 1852 8132 1858 8134
rect 1550 8123 1858 8132
rect 5550 8188 5858 8197
rect 5550 8186 5556 8188
rect 5612 8186 5636 8188
rect 5692 8186 5716 8188
rect 5772 8186 5796 8188
rect 5852 8186 5858 8188
rect 5612 8134 5614 8186
rect 5794 8134 5796 8186
rect 5550 8132 5556 8134
rect 5612 8132 5636 8134
rect 5692 8132 5716 8134
rect 5772 8132 5796 8134
rect 5852 8132 5858 8134
rect 5550 8123 5858 8132
rect 9550 8188 9858 8197
rect 9550 8186 9556 8188
rect 9612 8186 9636 8188
rect 9692 8186 9716 8188
rect 9772 8186 9796 8188
rect 9852 8186 9858 8188
rect 9612 8134 9614 8186
rect 9794 8134 9796 8186
rect 9550 8132 9556 8134
rect 9612 8132 9636 8134
rect 9692 8132 9716 8134
rect 9772 8132 9796 8134
rect 9852 8132 9858 8134
rect 9550 8123 9858 8132
rect 13550 8188 13858 8197
rect 13550 8186 13556 8188
rect 13612 8186 13636 8188
rect 13692 8186 13716 8188
rect 13772 8186 13796 8188
rect 13852 8186 13858 8188
rect 13612 8134 13614 8186
rect 13794 8134 13796 8186
rect 13550 8132 13556 8134
rect 13612 8132 13636 8134
rect 13692 8132 13716 8134
rect 13772 8132 13796 8134
rect 13852 8132 13858 8134
rect 13550 8123 13858 8132
rect 17550 8188 17858 8197
rect 17550 8186 17556 8188
rect 17612 8186 17636 8188
rect 17692 8186 17716 8188
rect 17772 8186 17796 8188
rect 17852 8186 17858 8188
rect 17612 8134 17614 8186
rect 17794 8134 17796 8186
rect 17550 8132 17556 8134
rect 17612 8132 17636 8134
rect 17692 8132 17716 8134
rect 17772 8132 17796 8134
rect 17852 8132 17858 8134
rect 17550 8123 17858 8132
rect 2210 7644 2518 7653
rect 2210 7642 2216 7644
rect 2272 7642 2296 7644
rect 2352 7642 2376 7644
rect 2432 7642 2456 7644
rect 2512 7642 2518 7644
rect 2272 7590 2274 7642
rect 2454 7590 2456 7642
rect 2210 7588 2216 7590
rect 2272 7588 2296 7590
rect 2352 7588 2376 7590
rect 2432 7588 2456 7590
rect 2512 7588 2518 7590
rect 2210 7579 2518 7588
rect 6210 7644 6518 7653
rect 6210 7642 6216 7644
rect 6272 7642 6296 7644
rect 6352 7642 6376 7644
rect 6432 7642 6456 7644
rect 6512 7642 6518 7644
rect 6272 7590 6274 7642
rect 6454 7590 6456 7642
rect 6210 7588 6216 7590
rect 6272 7588 6296 7590
rect 6352 7588 6376 7590
rect 6432 7588 6456 7590
rect 6512 7588 6518 7590
rect 6210 7579 6518 7588
rect 10210 7644 10518 7653
rect 10210 7642 10216 7644
rect 10272 7642 10296 7644
rect 10352 7642 10376 7644
rect 10432 7642 10456 7644
rect 10512 7642 10518 7644
rect 10272 7590 10274 7642
rect 10454 7590 10456 7642
rect 10210 7588 10216 7590
rect 10272 7588 10296 7590
rect 10352 7588 10376 7590
rect 10432 7588 10456 7590
rect 10512 7588 10518 7590
rect 10210 7579 10518 7588
rect 14210 7644 14518 7653
rect 14210 7642 14216 7644
rect 14272 7642 14296 7644
rect 14352 7642 14376 7644
rect 14432 7642 14456 7644
rect 14512 7642 14518 7644
rect 14272 7590 14274 7642
rect 14454 7590 14456 7642
rect 14210 7588 14216 7590
rect 14272 7588 14296 7590
rect 14352 7588 14376 7590
rect 14432 7588 14456 7590
rect 14512 7588 14518 7590
rect 14210 7579 14518 7588
rect 18210 7644 18518 7653
rect 18210 7642 18216 7644
rect 18272 7642 18296 7644
rect 18352 7642 18376 7644
rect 18432 7642 18456 7644
rect 18512 7642 18518 7644
rect 18272 7590 18274 7642
rect 18454 7590 18456 7642
rect 18210 7588 18216 7590
rect 18272 7588 18296 7590
rect 18352 7588 18376 7590
rect 18432 7588 18456 7590
rect 18512 7588 18518 7590
rect 18210 7579 18518 7588
rect 1550 7100 1858 7109
rect 1550 7098 1556 7100
rect 1612 7098 1636 7100
rect 1692 7098 1716 7100
rect 1772 7098 1796 7100
rect 1852 7098 1858 7100
rect 1612 7046 1614 7098
rect 1794 7046 1796 7098
rect 1550 7044 1556 7046
rect 1612 7044 1636 7046
rect 1692 7044 1716 7046
rect 1772 7044 1796 7046
rect 1852 7044 1858 7046
rect 1550 7035 1858 7044
rect 5550 7100 5858 7109
rect 5550 7098 5556 7100
rect 5612 7098 5636 7100
rect 5692 7098 5716 7100
rect 5772 7098 5796 7100
rect 5852 7098 5858 7100
rect 5612 7046 5614 7098
rect 5794 7046 5796 7098
rect 5550 7044 5556 7046
rect 5612 7044 5636 7046
rect 5692 7044 5716 7046
rect 5772 7044 5796 7046
rect 5852 7044 5858 7046
rect 5550 7035 5858 7044
rect 9550 7100 9858 7109
rect 9550 7098 9556 7100
rect 9612 7098 9636 7100
rect 9692 7098 9716 7100
rect 9772 7098 9796 7100
rect 9852 7098 9858 7100
rect 9612 7046 9614 7098
rect 9794 7046 9796 7098
rect 9550 7044 9556 7046
rect 9612 7044 9636 7046
rect 9692 7044 9716 7046
rect 9772 7044 9796 7046
rect 9852 7044 9858 7046
rect 9550 7035 9858 7044
rect 13550 7100 13858 7109
rect 13550 7098 13556 7100
rect 13612 7098 13636 7100
rect 13692 7098 13716 7100
rect 13772 7098 13796 7100
rect 13852 7098 13858 7100
rect 13612 7046 13614 7098
rect 13794 7046 13796 7098
rect 13550 7044 13556 7046
rect 13612 7044 13636 7046
rect 13692 7044 13716 7046
rect 13772 7044 13796 7046
rect 13852 7044 13858 7046
rect 13550 7035 13858 7044
rect 17550 7100 17858 7109
rect 17550 7098 17556 7100
rect 17612 7098 17636 7100
rect 17692 7098 17716 7100
rect 17772 7098 17796 7100
rect 17852 7098 17858 7100
rect 17612 7046 17614 7098
rect 17794 7046 17796 7098
rect 17550 7044 17556 7046
rect 17612 7044 17636 7046
rect 17692 7044 17716 7046
rect 17772 7044 17796 7046
rect 17852 7044 17858 7046
rect 17550 7035 17858 7044
rect 2210 6556 2518 6565
rect 2210 6554 2216 6556
rect 2272 6554 2296 6556
rect 2352 6554 2376 6556
rect 2432 6554 2456 6556
rect 2512 6554 2518 6556
rect 2272 6502 2274 6554
rect 2454 6502 2456 6554
rect 2210 6500 2216 6502
rect 2272 6500 2296 6502
rect 2352 6500 2376 6502
rect 2432 6500 2456 6502
rect 2512 6500 2518 6502
rect 2210 6491 2518 6500
rect 6210 6556 6518 6565
rect 6210 6554 6216 6556
rect 6272 6554 6296 6556
rect 6352 6554 6376 6556
rect 6432 6554 6456 6556
rect 6512 6554 6518 6556
rect 6272 6502 6274 6554
rect 6454 6502 6456 6554
rect 6210 6500 6216 6502
rect 6272 6500 6296 6502
rect 6352 6500 6376 6502
rect 6432 6500 6456 6502
rect 6512 6500 6518 6502
rect 6210 6491 6518 6500
rect 10210 6556 10518 6565
rect 10210 6554 10216 6556
rect 10272 6554 10296 6556
rect 10352 6554 10376 6556
rect 10432 6554 10456 6556
rect 10512 6554 10518 6556
rect 10272 6502 10274 6554
rect 10454 6502 10456 6554
rect 10210 6500 10216 6502
rect 10272 6500 10296 6502
rect 10352 6500 10376 6502
rect 10432 6500 10456 6502
rect 10512 6500 10518 6502
rect 10210 6491 10518 6500
rect 14210 6556 14518 6565
rect 14210 6554 14216 6556
rect 14272 6554 14296 6556
rect 14352 6554 14376 6556
rect 14432 6554 14456 6556
rect 14512 6554 14518 6556
rect 14272 6502 14274 6554
rect 14454 6502 14456 6554
rect 14210 6500 14216 6502
rect 14272 6500 14296 6502
rect 14352 6500 14376 6502
rect 14432 6500 14456 6502
rect 14512 6500 14518 6502
rect 14210 6491 14518 6500
rect 18210 6556 18518 6565
rect 18210 6554 18216 6556
rect 18272 6554 18296 6556
rect 18352 6554 18376 6556
rect 18432 6554 18456 6556
rect 18512 6554 18518 6556
rect 18272 6502 18274 6554
rect 18454 6502 18456 6554
rect 18210 6500 18216 6502
rect 18272 6500 18296 6502
rect 18352 6500 18376 6502
rect 18432 6500 18456 6502
rect 18512 6500 18518 6502
rect 18210 6491 18518 6500
rect 1550 6012 1858 6021
rect 1550 6010 1556 6012
rect 1612 6010 1636 6012
rect 1692 6010 1716 6012
rect 1772 6010 1796 6012
rect 1852 6010 1858 6012
rect 1612 5958 1614 6010
rect 1794 5958 1796 6010
rect 1550 5956 1556 5958
rect 1612 5956 1636 5958
rect 1692 5956 1716 5958
rect 1772 5956 1796 5958
rect 1852 5956 1858 5958
rect 1550 5947 1858 5956
rect 5550 6012 5858 6021
rect 5550 6010 5556 6012
rect 5612 6010 5636 6012
rect 5692 6010 5716 6012
rect 5772 6010 5796 6012
rect 5852 6010 5858 6012
rect 5612 5958 5614 6010
rect 5794 5958 5796 6010
rect 5550 5956 5556 5958
rect 5612 5956 5636 5958
rect 5692 5956 5716 5958
rect 5772 5956 5796 5958
rect 5852 5956 5858 5958
rect 5550 5947 5858 5956
rect 9550 6012 9858 6021
rect 9550 6010 9556 6012
rect 9612 6010 9636 6012
rect 9692 6010 9716 6012
rect 9772 6010 9796 6012
rect 9852 6010 9858 6012
rect 9612 5958 9614 6010
rect 9794 5958 9796 6010
rect 9550 5956 9556 5958
rect 9612 5956 9636 5958
rect 9692 5956 9716 5958
rect 9772 5956 9796 5958
rect 9852 5956 9858 5958
rect 9550 5947 9858 5956
rect 13550 6012 13858 6021
rect 13550 6010 13556 6012
rect 13612 6010 13636 6012
rect 13692 6010 13716 6012
rect 13772 6010 13796 6012
rect 13852 6010 13858 6012
rect 13612 5958 13614 6010
rect 13794 5958 13796 6010
rect 13550 5956 13556 5958
rect 13612 5956 13636 5958
rect 13692 5956 13716 5958
rect 13772 5956 13796 5958
rect 13852 5956 13858 5958
rect 13550 5947 13858 5956
rect 17550 6012 17858 6021
rect 17550 6010 17556 6012
rect 17612 6010 17636 6012
rect 17692 6010 17716 6012
rect 17772 6010 17796 6012
rect 17852 6010 17858 6012
rect 17612 5958 17614 6010
rect 17794 5958 17796 6010
rect 17550 5956 17556 5958
rect 17612 5956 17636 5958
rect 17692 5956 17716 5958
rect 17772 5956 17796 5958
rect 17852 5956 17858 5958
rect 17550 5947 17858 5956
rect 2210 5468 2518 5477
rect 2210 5466 2216 5468
rect 2272 5466 2296 5468
rect 2352 5466 2376 5468
rect 2432 5466 2456 5468
rect 2512 5466 2518 5468
rect 2272 5414 2274 5466
rect 2454 5414 2456 5466
rect 2210 5412 2216 5414
rect 2272 5412 2296 5414
rect 2352 5412 2376 5414
rect 2432 5412 2456 5414
rect 2512 5412 2518 5414
rect 2210 5403 2518 5412
rect 6210 5468 6518 5477
rect 6210 5466 6216 5468
rect 6272 5466 6296 5468
rect 6352 5466 6376 5468
rect 6432 5466 6456 5468
rect 6512 5466 6518 5468
rect 6272 5414 6274 5466
rect 6454 5414 6456 5466
rect 6210 5412 6216 5414
rect 6272 5412 6296 5414
rect 6352 5412 6376 5414
rect 6432 5412 6456 5414
rect 6512 5412 6518 5414
rect 6210 5403 6518 5412
rect 10210 5468 10518 5477
rect 10210 5466 10216 5468
rect 10272 5466 10296 5468
rect 10352 5466 10376 5468
rect 10432 5466 10456 5468
rect 10512 5466 10518 5468
rect 10272 5414 10274 5466
rect 10454 5414 10456 5466
rect 10210 5412 10216 5414
rect 10272 5412 10296 5414
rect 10352 5412 10376 5414
rect 10432 5412 10456 5414
rect 10512 5412 10518 5414
rect 10210 5403 10518 5412
rect 14210 5468 14518 5477
rect 14210 5466 14216 5468
rect 14272 5466 14296 5468
rect 14352 5466 14376 5468
rect 14432 5466 14456 5468
rect 14512 5466 14518 5468
rect 14272 5414 14274 5466
rect 14454 5414 14456 5466
rect 14210 5412 14216 5414
rect 14272 5412 14296 5414
rect 14352 5412 14376 5414
rect 14432 5412 14456 5414
rect 14512 5412 14518 5414
rect 14210 5403 14518 5412
rect 18210 5468 18518 5477
rect 18210 5466 18216 5468
rect 18272 5466 18296 5468
rect 18352 5466 18376 5468
rect 18432 5466 18456 5468
rect 18512 5466 18518 5468
rect 18272 5414 18274 5466
rect 18454 5414 18456 5466
rect 18210 5412 18216 5414
rect 18272 5412 18296 5414
rect 18352 5412 18376 5414
rect 18432 5412 18456 5414
rect 18512 5412 18518 5414
rect 18210 5403 18518 5412
rect 1550 4924 1858 4933
rect 1550 4922 1556 4924
rect 1612 4922 1636 4924
rect 1692 4922 1716 4924
rect 1772 4922 1796 4924
rect 1852 4922 1858 4924
rect 1612 4870 1614 4922
rect 1794 4870 1796 4922
rect 1550 4868 1556 4870
rect 1612 4868 1636 4870
rect 1692 4868 1716 4870
rect 1772 4868 1796 4870
rect 1852 4868 1858 4870
rect 1550 4859 1858 4868
rect 5550 4924 5858 4933
rect 5550 4922 5556 4924
rect 5612 4922 5636 4924
rect 5692 4922 5716 4924
rect 5772 4922 5796 4924
rect 5852 4922 5858 4924
rect 5612 4870 5614 4922
rect 5794 4870 5796 4922
rect 5550 4868 5556 4870
rect 5612 4868 5636 4870
rect 5692 4868 5716 4870
rect 5772 4868 5796 4870
rect 5852 4868 5858 4870
rect 5550 4859 5858 4868
rect 9550 4924 9858 4933
rect 9550 4922 9556 4924
rect 9612 4922 9636 4924
rect 9692 4922 9716 4924
rect 9772 4922 9796 4924
rect 9852 4922 9858 4924
rect 9612 4870 9614 4922
rect 9794 4870 9796 4922
rect 9550 4868 9556 4870
rect 9612 4868 9636 4870
rect 9692 4868 9716 4870
rect 9772 4868 9796 4870
rect 9852 4868 9858 4870
rect 9550 4859 9858 4868
rect 13550 4924 13858 4933
rect 13550 4922 13556 4924
rect 13612 4922 13636 4924
rect 13692 4922 13716 4924
rect 13772 4922 13796 4924
rect 13852 4922 13858 4924
rect 13612 4870 13614 4922
rect 13794 4870 13796 4922
rect 13550 4868 13556 4870
rect 13612 4868 13636 4870
rect 13692 4868 13716 4870
rect 13772 4868 13796 4870
rect 13852 4868 13858 4870
rect 13550 4859 13858 4868
rect 17550 4924 17858 4933
rect 17550 4922 17556 4924
rect 17612 4922 17636 4924
rect 17692 4922 17716 4924
rect 17772 4922 17796 4924
rect 17852 4922 17858 4924
rect 17612 4870 17614 4922
rect 17794 4870 17796 4922
rect 17550 4868 17556 4870
rect 17612 4868 17636 4870
rect 17692 4868 17716 4870
rect 17772 4868 17796 4870
rect 17852 4868 17858 4870
rect 17550 4859 17858 4868
rect 2210 4380 2518 4389
rect 2210 4378 2216 4380
rect 2272 4378 2296 4380
rect 2352 4378 2376 4380
rect 2432 4378 2456 4380
rect 2512 4378 2518 4380
rect 2272 4326 2274 4378
rect 2454 4326 2456 4378
rect 2210 4324 2216 4326
rect 2272 4324 2296 4326
rect 2352 4324 2376 4326
rect 2432 4324 2456 4326
rect 2512 4324 2518 4326
rect 2210 4315 2518 4324
rect 6210 4380 6518 4389
rect 6210 4378 6216 4380
rect 6272 4378 6296 4380
rect 6352 4378 6376 4380
rect 6432 4378 6456 4380
rect 6512 4378 6518 4380
rect 6272 4326 6274 4378
rect 6454 4326 6456 4378
rect 6210 4324 6216 4326
rect 6272 4324 6296 4326
rect 6352 4324 6376 4326
rect 6432 4324 6456 4326
rect 6512 4324 6518 4326
rect 6210 4315 6518 4324
rect 10210 4380 10518 4389
rect 10210 4378 10216 4380
rect 10272 4378 10296 4380
rect 10352 4378 10376 4380
rect 10432 4378 10456 4380
rect 10512 4378 10518 4380
rect 10272 4326 10274 4378
rect 10454 4326 10456 4378
rect 10210 4324 10216 4326
rect 10272 4324 10296 4326
rect 10352 4324 10376 4326
rect 10432 4324 10456 4326
rect 10512 4324 10518 4326
rect 10210 4315 10518 4324
rect 14210 4380 14518 4389
rect 14210 4378 14216 4380
rect 14272 4378 14296 4380
rect 14352 4378 14376 4380
rect 14432 4378 14456 4380
rect 14512 4378 14518 4380
rect 14272 4326 14274 4378
rect 14454 4326 14456 4378
rect 14210 4324 14216 4326
rect 14272 4324 14296 4326
rect 14352 4324 14376 4326
rect 14432 4324 14456 4326
rect 14512 4324 14518 4326
rect 14210 4315 14518 4324
rect 18210 4380 18518 4389
rect 18210 4378 18216 4380
rect 18272 4378 18296 4380
rect 18352 4378 18376 4380
rect 18432 4378 18456 4380
rect 18512 4378 18518 4380
rect 18272 4326 18274 4378
rect 18454 4326 18456 4378
rect 18210 4324 18216 4326
rect 18272 4324 18296 4326
rect 18352 4324 18376 4326
rect 18432 4324 18456 4326
rect 18512 4324 18518 4326
rect 18210 4315 18518 4324
rect 1550 3836 1858 3845
rect 1550 3834 1556 3836
rect 1612 3834 1636 3836
rect 1692 3834 1716 3836
rect 1772 3834 1796 3836
rect 1852 3834 1858 3836
rect 1612 3782 1614 3834
rect 1794 3782 1796 3834
rect 1550 3780 1556 3782
rect 1612 3780 1636 3782
rect 1692 3780 1716 3782
rect 1772 3780 1796 3782
rect 1852 3780 1858 3782
rect 1550 3771 1858 3780
rect 5550 3836 5858 3845
rect 5550 3834 5556 3836
rect 5612 3834 5636 3836
rect 5692 3834 5716 3836
rect 5772 3834 5796 3836
rect 5852 3834 5858 3836
rect 5612 3782 5614 3834
rect 5794 3782 5796 3834
rect 5550 3780 5556 3782
rect 5612 3780 5636 3782
rect 5692 3780 5716 3782
rect 5772 3780 5796 3782
rect 5852 3780 5858 3782
rect 5550 3771 5858 3780
rect 9550 3836 9858 3845
rect 9550 3834 9556 3836
rect 9612 3834 9636 3836
rect 9692 3834 9716 3836
rect 9772 3834 9796 3836
rect 9852 3834 9858 3836
rect 9612 3782 9614 3834
rect 9794 3782 9796 3834
rect 9550 3780 9556 3782
rect 9612 3780 9636 3782
rect 9692 3780 9716 3782
rect 9772 3780 9796 3782
rect 9852 3780 9858 3782
rect 9550 3771 9858 3780
rect 13550 3836 13858 3845
rect 13550 3834 13556 3836
rect 13612 3834 13636 3836
rect 13692 3834 13716 3836
rect 13772 3834 13796 3836
rect 13852 3834 13858 3836
rect 13612 3782 13614 3834
rect 13794 3782 13796 3834
rect 13550 3780 13556 3782
rect 13612 3780 13636 3782
rect 13692 3780 13716 3782
rect 13772 3780 13796 3782
rect 13852 3780 13858 3782
rect 13550 3771 13858 3780
rect 17550 3836 17858 3845
rect 17550 3834 17556 3836
rect 17612 3834 17636 3836
rect 17692 3834 17716 3836
rect 17772 3834 17796 3836
rect 17852 3834 17858 3836
rect 17612 3782 17614 3834
rect 17794 3782 17796 3834
rect 17550 3780 17556 3782
rect 17612 3780 17636 3782
rect 17692 3780 17716 3782
rect 17772 3780 17796 3782
rect 17852 3780 17858 3782
rect 17550 3771 17858 3780
rect 2210 3292 2518 3301
rect 2210 3290 2216 3292
rect 2272 3290 2296 3292
rect 2352 3290 2376 3292
rect 2432 3290 2456 3292
rect 2512 3290 2518 3292
rect 2272 3238 2274 3290
rect 2454 3238 2456 3290
rect 2210 3236 2216 3238
rect 2272 3236 2296 3238
rect 2352 3236 2376 3238
rect 2432 3236 2456 3238
rect 2512 3236 2518 3238
rect 2210 3227 2518 3236
rect 6210 3292 6518 3301
rect 6210 3290 6216 3292
rect 6272 3290 6296 3292
rect 6352 3290 6376 3292
rect 6432 3290 6456 3292
rect 6512 3290 6518 3292
rect 6272 3238 6274 3290
rect 6454 3238 6456 3290
rect 6210 3236 6216 3238
rect 6272 3236 6296 3238
rect 6352 3236 6376 3238
rect 6432 3236 6456 3238
rect 6512 3236 6518 3238
rect 6210 3227 6518 3236
rect 10210 3292 10518 3301
rect 10210 3290 10216 3292
rect 10272 3290 10296 3292
rect 10352 3290 10376 3292
rect 10432 3290 10456 3292
rect 10512 3290 10518 3292
rect 10272 3238 10274 3290
rect 10454 3238 10456 3290
rect 10210 3236 10216 3238
rect 10272 3236 10296 3238
rect 10352 3236 10376 3238
rect 10432 3236 10456 3238
rect 10512 3236 10518 3238
rect 10210 3227 10518 3236
rect 14210 3292 14518 3301
rect 14210 3290 14216 3292
rect 14272 3290 14296 3292
rect 14352 3290 14376 3292
rect 14432 3290 14456 3292
rect 14512 3290 14518 3292
rect 14272 3238 14274 3290
rect 14454 3238 14456 3290
rect 14210 3236 14216 3238
rect 14272 3236 14296 3238
rect 14352 3236 14376 3238
rect 14432 3236 14456 3238
rect 14512 3236 14518 3238
rect 14210 3227 14518 3236
rect 18210 3292 18518 3301
rect 18210 3290 18216 3292
rect 18272 3290 18296 3292
rect 18352 3290 18376 3292
rect 18432 3290 18456 3292
rect 18512 3290 18518 3292
rect 18272 3238 18274 3290
rect 18454 3238 18456 3290
rect 18210 3236 18216 3238
rect 18272 3236 18296 3238
rect 18352 3236 18376 3238
rect 18432 3236 18456 3238
rect 18512 3236 18518 3238
rect 18210 3227 18518 3236
rect 1550 2748 1858 2757
rect 1550 2746 1556 2748
rect 1612 2746 1636 2748
rect 1692 2746 1716 2748
rect 1772 2746 1796 2748
rect 1852 2746 1858 2748
rect 1612 2694 1614 2746
rect 1794 2694 1796 2746
rect 1550 2692 1556 2694
rect 1612 2692 1636 2694
rect 1692 2692 1716 2694
rect 1772 2692 1796 2694
rect 1852 2692 1858 2694
rect 1550 2683 1858 2692
rect 5550 2748 5858 2757
rect 5550 2746 5556 2748
rect 5612 2746 5636 2748
rect 5692 2746 5716 2748
rect 5772 2746 5796 2748
rect 5852 2746 5858 2748
rect 5612 2694 5614 2746
rect 5794 2694 5796 2746
rect 5550 2692 5556 2694
rect 5612 2692 5636 2694
rect 5692 2692 5716 2694
rect 5772 2692 5796 2694
rect 5852 2692 5858 2694
rect 5550 2683 5858 2692
rect 9550 2748 9858 2757
rect 9550 2746 9556 2748
rect 9612 2746 9636 2748
rect 9692 2746 9716 2748
rect 9772 2746 9796 2748
rect 9852 2746 9858 2748
rect 9612 2694 9614 2746
rect 9794 2694 9796 2746
rect 9550 2692 9556 2694
rect 9612 2692 9636 2694
rect 9692 2692 9716 2694
rect 9772 2692 9796 2694
rect 9852 2692 9858 2694
rect 9550 2683 9858 2692
rect 13550 2748 13858 2757
rect 13550 2746 13556 2748
rect 13612 2746 13636 2748
rect 13692 2746 13716 2748
rect 13772 2746 13796 2748
rect 13852 2746 13858 2748
rect 13612 2694 13614 2746
rect 13794 2694 13796 2746
rect 13550 2692 13556 2694
rect 13612 2692 13636 2694
rect 13692 2692 13716 2694
rect 13772 2692 13796 2694
rect 13852 2692 13858 2694
rect 13550 2683 13858 2692
rect 17550 2748 17858 2757
rect 17550 2746 17556 2748
rect 17612 2746 17636 2748
rect 17692 2746 17716 2748
rect 17772 2746 17796 2748
rect 17852 2746 17858 2748
rect 17612 2694 17614 2746
rect 17794 2694 17796 2746
rect 17550 2692 17556 2694
rect 17612 2692 17636 2694
rect 17692 2692 17716 2694
rect 17772 2692 17796 2694
rect 17852 2692 17858 2694
rect 17550 2683 17858 2692
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 2210 2204 2518 2213
rect 2210 2202 2216 2204
rect 2272 2202 2296 2204
rect 2352 2202 2376 2204
rect 2432 2202 2456 2204
rect 2512 2202 2518 2204
rect 2272 2150 2274 2202
rect 2454 2150 2456 2202
rect 2210 2148 2216 2150
rect 2272 2148 2296 2150
rect 2352 2148 2376 2150
rect 2432 2148 2456 2150
rect 2512 2148 2518 2150
rect 2210 2139 2518 2148
rect 6210 2204 6518 2213
rect 6210 2202 6216 2204
rect 6272 2202 6296 2204
rect 6352 2202 6376 2204
rect 6432 2202 6456 2204
rect 6512 2202 6518 2204
rect 6272 2150 6274 2202
rect 6454 2150 6456 2202
rect 6210 2148 6216 2150
rect 6272 2148 6296 2150
rect 6352 2148 6376 2150
rect 6432 2148 6456 2150
rect 6512 2148 6518 2150
rect 6210 2139 6518 2148
rect 9692 800 9720 2382
rect 10152 1306 10180 2382
rect 10210 2204 10518 2213
rect 10210 2202 10216 2204
rect 10272 2202 10296 2204
rect 10352 2202 10376 2204
rect 10432 2202 10456 2204
rect 10512 2202 10518 2204
rect 10272 2150 10274 2202
rect 10454 2150 10456 2202
rect 10210 2148 10216 2150
rect 10272 2148 10296 2150
rect 10352 2148 10376 2150
rect 10432 2148 10456 2150
rect 10512 2148 10518 2150
rect 10210 2139 10518 2148
rect 14210 2204 14518 2213
rect 14210 2202 14216 2204
rect 14272 2202 14296 2204
rect 14352 2202 14376 2204
rect 14432 2202 14456 2204
rect 14512 2202 14518 2204
rect 14272 2150 14274 2202
rect 14454 2150 14456 2202
rect 14210 2148 14216 2150
rect 14272 2148 14296 2150
rect 14352 2148 14376 2150
rect 14432 2148 14456 2150
rect 14512 2148 14518 2150
rect 14210 2139 14518 2148
rect 18210 2204 18518 2213
rect 18210 2202 18216 2204
rect 18272 2202 18296 2204
rect 18352 2202 18376 2204
rect 18432 2202 18456 2204
rect 18512 2202 18518 2204
rect 18272 2150 18274 2202
rect 18454 2150 18456 2202
rect 18210 2148 18216 2150
rect 18272 2148 18296 2150
rect 18352 2148 18376 2150
rect 18432 2148 18456 2150
rect 18512 2148 18518 2150
rect 18210 2139 18518 2148
rect 10152 1278 10364 1306
rect 10336 800 10364 1278
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 9678 0 9734 800
rect 10322 0 10378 800
<< via2 >>
rect 2216 17434 2272 17436
rect 2296 17434 2352 17436
rect 2376 17434 2432 17436
rect 2456 17434 2512 17436
rect 2216 17382 2262 17434
rect 2262 17382 2272 17434
rect 2296 17382 2326 17434
rect 2326 17382 2338 17434
rect 2338 17382 2352 17434
rect 2376 17382 2390 17434
rect 2390 17382 2402 17434
rect 2402 17382 2432 17434
rect 2456 17382 2466 17434
rect 2466 17382 2512 17434
rect 2216 17380 2272 17382
rect 2296 17380 2352 17382
rect 2376 17380 2432 17382
rect 2456 17380 2512 17382
rect 6216 17434 6272 17436
rect 6296 17434 6352 17436
rect 6376 17434 6432 17436
rect 6456 17434 6512 17436
rect 6216 17382 6262 17434
rect 6262 17382 6272 17434
rect 6296 17382 6326 17434
rect 6326 17382 6338 17434
rect 6338 17382 6352 17434
rect 6376 17382 6390 17434
rect 6390 17382 6402 17434
rect 6402 17382 6432 17434
rect 6456 17382 6466 17434
rect 6466 17382 6512 17434
rect 6216 17380 6272 17382
rect 6296 17380 6352 17382
rect 6376 17380 6432 17382
rect 6456 17380 6512 17382
rect 10216 17434 10272 17436
rect 10296 17434 10352 17436
rect 10376 17434 10432 17436
rect 10456 17434 10512 17436
rect 10216 17382 10262 17434
rect 10262 17382 10272 17434
rect 10296 17382 10326 17434
rect 10326 17382 10338 17434
rect 10338 17382 10352 17434
rect 10376 17382 10390 17434
rect 10390 17382 10402 17434
rect 10402 17382 10432 17434
rect 10456 17382 10466 17434
rect 10466 17382 10512 17434
rect 10216 17380 10272 17382
rect 10296 17380 10352 17382
rect 10376 17380 10432 17382
rect 10456 17380 10512 17382
rect 14216 17434 14272 17436
rect 14296 17434 14352 17436
rect 14376 17434 14432 17436
rect 14456 17434 14512 17436
rect 14216 17382 14262 17434
rect 14262 17382 14272 17434
rect 14296 17382 14326 17434
rect 14326 17382 14338 17434
rect 14338 17382 14352 17434
rect 14376 17382 14390 17434
rect 14390 17382 14402 17434
rect 14402 17382 14432 17434
rect 14456 17382 14466 17434
rect 14466 17382 14512 17434
rect 14216 17380 14272 17382
rect 14296 17380 14352 17382
rect 14376 17380 14432 17382
rect 14456 17380 14512 17382
rect 18216 17434 18272 17436
rect 18296 17434 18352 17436
rect 18376 17434 18432 17436
rect 18456 17434 18512 17436
rect 18216 17382 18262 17434
rect 18262 17382 18272 17434
rect 18296 17382 18326 17434
rect 18326 17382 18338 17434
rect 18338 17382 18352 17434
rect 18376 17382 18390 17434
rect 18390 17382 18402 17434
rect 18402 17382 18432 17434
rect 18456 17382 18466 17434
rect 18466 17382 18512 17434
rect 18216 17380 18272 17382
rect 18296 17380 18352 17382
rect 18376 17380 18432 17382
rect 18456 17380 18512 17382
rect 1556 16890 1612 16892
rect 1636 16890 1692 16892
rect 1716 16890 1772 16892
rect 1796 16890 1852 16892
rect 1556 16838 1602 16890
rect 1602 16838 1612 16890
rect 1636 16838 1666 16890
rect 1666 16838 1678 16890
rect 1678 16838 1692 16890
rect 1716 16838 1730 16890
rect 1730 16838 1742 16890
rect 1742 16838 1772 16890
rect 1796 16838 1806 16890
rect 1806 16838 1852 16890
rect 1556 16836 1612 16838
rect 1636 16836 1692 16838
rect 1716 16836 1772 16838
rect 1796 16836 1852 16838
rect 5556 16890 5612 16892
rect 5636 16890 5692 16892
rect 5716 16890 5772 16892
rect 5796 16890 5852 16892
rect 5556 16838 5602 16890
rect 5602 16838 5612 16890
rect 5636 16838 5666 16890
rect 5666 16838 5678 16890
rect 5678 16838 5692 16890
rect 5716 16838 5730 16890
rect 5730 16838 5742 16890
rect 5742 16838 5772 16890
rect 5796 16838 5806 16890
rect 5806 16838 5852 16890
rect 5556 16836 5612 16838
rect 5636 16836 5692 16838
rect 5716 16836 5772 16838
rect 5796 16836 5852 16838
rect 9556 16890 9612 16892
rect 9636 16890 9692 16892
rect 9716 16890 9772 16892
rect 9796 16890 9852 16892
rect 9556 16838 9602 16890
rect 9602 16838 9612 16890
rect 9636 16838 9666 16890
rect 9666 16838 9678 16890
rect 9678 16838 9692 16890
rect 9716 16838 9730 16890
rect 9730 16838 9742 16890
rect 9742 16838 9772 16890
rect 9796 16838 9806 16890
rect 9806 16838 9852 16890
rect 9556 16836 9612 16838
rect 9636 16836 9692 16838
rect 9716 16836 9772 16838
rect 9796 16836 9852 16838
rect 13556 16890 13612 16892
rect 13636 16890 13692 16892
rect 13716 16890 13772 16892
rect 13796 16890 13852 16892
rect 13556 16838 13602 16890
rect 13602 16838 13612 16890
rect 13636 16838 13666 16890
rect 13666 16838 13678 16890
rect 13678 16838 13692 16890
rect 13716 16838 13730 16890
rect 13730 16838 13742 16890
rect 13742 16838 13772 16890
rect 13796 16838 13806 16890
rect 13806 16838 13852 16890
rect 13556 16836 13612 16838
rect 13636 16836 13692 16838
rect 13716 16836 13772 16838
rect 13796 16836 13852 16838
rect 17556 16890 17612 16892
rect 17636 16890 17692 16892
rect 17716 16890 17772 16892
rect 17796 16890 17852 16892
rect 17556 16838 17602 16890
rect 17602 16838 17612 16890
rect 17636 16838 17666 16890
rect 17666 16838 17678 16890
rect 17678 16838 17692 16890
rect 17716 16838 17730 16890
rect 17730 16838 17742 16890
rect 17742 16838 17772 16890
rect 17796 16838 17806 16890
rect 17806 16838 17852 16890
rect 17556 16836 17612 16838
rect 17636 16836 17692 16838
rect 17716 16836 17772 16838
rect 17796 16836 17852 16838
rect 2216 16346 2272 16348
rect 2296 16346 2352 16348
rect 2376 16346 2432 16348
rect 2456 16346 2512 16348
rect 2216 16294 2262 16346
rect 2262 16294 2272 16346
rect 2296 16294 2326 16346
rect 2326 16294 2338 16346
rect 2338 16294 2352 16346
rect 2376 16294 2390 16346
rect 2390 16294 2402 16346
rect 2402 16294 2432 16346
rect 2456 16294 2466 16346
rect 2466 16294 2512 16346
rect 2216 16292 2272 16294
rect 2296 16292 2352 16294
rect 2376 16292 2432 16294
rect 2456 16292 2512 16294
rect 6216 16346 6272 16348
rect 6296 16346 6352 16348
rect 6376 16346 6432 16348
rect 6456 16346 6512 16348
rect 6216 16294 6262 16346
rect 6262 16294 6272 16346
rect 6296 16294 6326 16346
rect 6326 16294 6338 16346
rect 6338 16294 6352 16346
rect 6376 16294 6390 16346
rect 6390 16294 6402 16346
rect 6402 16294 6432 16346
rect 6456 16294 6466 16346
rect 6466 16294 6512 16346
rect 6216 16292 6272 16294
rect 6296 16292 6352 16294
rect 6376 16292 6432 16294
rect 6456 16292 6512 16294
rect 10216 16346 10272 16348
rect 10296 16346 10352 16348
rect 10376 16346 10432 16348
rect 10456 16346 10512 16348
rect 10216 16294 10262 16346
rect 10262 16294 10272 16346
rect 10296 16294 10326 16346
rect 10326 16294 10338 16346
rect 10338 16294 10352 16346
rect 10376 16294 10390 16346
rect 10390 16294 10402 16346
rect 10402 16294 10432 16346
rect 10456 16294 10466 16346
rect 10466 16294 10512 16346
rect 10216 16292 10272 16294
rect 10296 16292 10352 16294
rect 10376 16292 10432 16294
rect 10456 16292 10512 16294
rect 14216 16346 14272 16348
rect 14296 16346 14352 16348
rect 14376 16346 14432 16348
rect 14456 16346 14512 16348
rect 14216 16294 14262 16346
rect 14262 16294 14272 16346
rect 14296 16294 14326 16346
rect 14326 16294 14338 16346
rect 14338 16294 14352 16346
rect 14376 16294 14390 16346
rect 14390 16294 14402 16346
rect 14402 16294 14432 16346
rect 14456 16294 14466 16346
rect 14466 16294 14512 16346
rect 14216 16292 14272 16294
rect 14296 16292 14352 16294
rect 14376 16292 14432 16294
rect 14456 16292 14512 16294
rect 18216 16346 18272 16348
rect 18296 16346 18352 16348
rect 18376 16346 18432 16348
rect 18456 16346 18512 16348
rect 18216 16294 18262 16346
rect 18262 16294 18272 16346
rect 18296 16294 18326 16346
rect 18326 16294 18338 16346
rect 18338 16294 18352 16346
rect 18376 16294 18390 16346
rect 18390 16294 18402 16346
rect 18402 16294 18432 16346
rect 18456 16294 18466 16346
rect 18466 16294 18512 16346
rect 18216 16292 18272 16294
rect 18296 16292 18352 16294
rect 18376 16292 18432 16294
rect 18456 16292 18512 16294
rect 1556 15802 1612 15804
rect 1636 15802 1692 15804
rect 1716 15802 1772 15804
rect 1796 15802 1852 15804
rect 1556 15750 1602 15802
rect 1602 15750 1612 15802
rect 1636 15750 1666 15802
rect 1666 15750 1678 15802
rect 1678 15750 1692 15802
rect 1716 15750 1730 15802
rect 1730 15750 1742 15802
rect 1742 15750 1772 15802
rect 1796 15750 1806 15802
rect 1806 15750 1852 15802
rect 1556 15748 1612 15750
rect 1636 15748 1692 15750
rect 1716 15748 1772 15750
rect 1796 15748 1852 15750
rect 5556 15802 5612 15804
rect 5636 15802 5692 15804
rect 5716 15802 5772 15804
rect 5796 15802 5852 15804
rect 5556 15750 5602 15802
rect 5602 15750 5612 15802
rect 5636 15750 5666 15802
rect 5666 15750 5678 15802
rect 5678 15750 5692 15802
rect 5716 15750 5730 15802
rect 5730 15750 5742 15802
rect 5742 15750 5772 15802
rect 5796 15750 5806 15802
rect 5806 15750 5852 15802
rect 5556 15748 5612 15750
rect 5636 15748 5692 15750
rect 5716 15748 5772 15750
rect 5796 15748 5852 15750
rect 9556 15802 9612 15804
rect 9636 15802 9692 15804
rect 9716 15802 9772 15804
rect 9796 15802 9852 15804
rect 9556 15750 9602 15802
rect 9602 15750 9612 15802
rect 9636 15750 9666 15802
rect 9666 15750 9678 15802
rect 9678 15750 9692 15802
rect 9716 15750 9730 15802
rect 9730 15750 9742 15802
rect 9742 15750 9772 15802
rect 9796 15750 9806 15802
rect 9806 15750 9852 15802
rect 9556 15748 9612 15750
rect 9636 15748 9692 15750
rect 9716 15748 9772 15750
rect 9796 15748 9852 15750
rect 13556 15802 13612 15804
rect 13636 15802 13692 15804
rect 13716 15802 13772 15804
rect 13796 15802 13852 15804
rect 13556 15750 13602 15802
rect 13602 15750 13612 15802
rect 13636 15750 13666 15802
rect 13666 15750 13678 15802
rect 13678 15750 13692 15802
rect 13716 15750 13730 15802
rect 13730 15750 13742 15802
rect 13742 15750 13772 15802
rect 13796 15750 13806 15802
rect 13806 15750 13852 15802
rect 13556 15748 13612 15750
rect 13636 15748 13692 15750
rect 13716 15748 13772 15750
rect 13796 15748 13852 15750
rect 17556 15802 17612 15804
rect 17636 15802 17692 15804
rect 17716 15802 17772 15804
rect 17796 15802 17852 15804
rect 17556 15750 17602 15802
rect 17602 15750 17612 15802
rect 17636 15750 17666 15802
rect 17666 15750 17678 15802
rect 17678 15750 17692 15802
rect 17716 15750 17730 15802
rect 17730 15750 17742 15802
rect 17742 15750 17772 15802
rect 17796 15750 17806 15802
rect 17806 15750 17852 15802
rect 17556 15748 17612 15750
rect 17636 15748 17692 15750
rect 17716 15748 17772 15750
rect 17796 15748 17852 15750
rect 2216 15258 2272 15260
rect 2296 15258 2352 15260
rect 2376 15258 2432 15260
rect 2456 15258 2512 15260
rect 2216 15206 2262 15258
rect 2262 15206 2272 15258
rect 2296 15206 2326 15258
rect 2326 15206 2338 15258
rect 2338 15206 2352 15258
rect 2376 15206 2390 15258
rect 2390 15206 2402 15258
rect 2402 15206 2432 15258
rect 2456 15206 2466 15258
rect 2466 15206 2512 15258
rect 2216 15204 2272 15206
rect 2296 15204 2352 15206
rect 2376 15204 2432 15206
rect 2456 15204 2512 15206
rect 6216 15258 6272 15260
rect 6296 15258 6352 15260
rect 6376 15258 6432 15260
rect 6456 15258 6512 15260
rect 6216 15206 6262 15258
rect 6262 15206 6272 15258
rect 6296 15206 6326 15258
rect 6326 15206 6338 15258
rect 6338 15206 6352 15258
rect 6376 15206 6390 15258
rect 6390 15206 6402 15258
rect 6402 15206 6432 15258
rect 6456 15206 6466 15258
rect 6466 15206 6512 15258
rect 6216 15204 6272 15206
rect 6296 15204 6352 15206
rect 6376 15204 6432 15206
rect 6456 15204 6512 15206
rect 10216 15258 10272 15260
rect 10296 15258 10352 15260
rect 10376 15258 10432 15260
rect 10456 15258 10512 15260
rect 10216 15206 10262 15258
rect 10262 15206 10272 15258
rect 10296 15206 10326 15258
rect 10326 15206 10338 15258
rect 10338 15206 10352 15258
rect 10376 15206 10390 15258
rect 10390 15206 10402 15258
rect 10402 15206 10432 15258
rect 10456 15206 10466 15258
rect 10466 15206 10512 15258
rect 10216 15204 10272 15206
rect 10296 15204 10352 15206
rect 10376 15204 10432 15206
rect 10456 15204 10512 15206
rect 14216 15258 14272 15260
rect 14296 15258 14352 15260
rect 14376 15258 14432 15260
rect 14456 15258 14512 15260
rect 14216 15206 14262 15258
rect 14262 15206 14272 15258
rect 14296 15206 14326 15258
rect 14326 15206 14338 15258
rect 14338 15206 14352 15258
rect 14376 15206 14390 15258
rect 14390 15206 14402 15258
rect 14402 15206 14432 15258
rect 14456 15206 14466 15258
rect 14466 15206 14512 15258
rect 14216 15204 14272 15206
rect 14296 15204 14352 15206
rect 14376 15204 14432 15206
rect 14456 15204 14512 15206
rect 18216 15258 18272 15260
rect 18296 15258 18352 15260
rect 18376 15258 18432 15260
rect 18456 15258 18512 15260
rect 18216 15206 18262 15258
rect 18262 15206 18272 15258
rect 18296 15206 18326 15258
rect 18326 15206 18338 15258
rect 18338 15206 18352 15258
rect 18376 15206 18390 15258
rect 18390 15206 18402 15258
rect 18402 15206 18432 15258
rect 18456 15206 18466 15258
rect 18466 15206 18512 15258
rect 18216 15204 18272 15206
rect 18296 15204 18352 15206
rect 18376 15204 18432 15206
rect 18456 15204 18512 15206
rect 1556 14714 1612 14716
rect 1636 14714 1692 14716
rect 1716 14714 1772 14716
rect 1796 14714 1852 14716
rect 1556 14662 1602 14714
rect 1602 14662 1612 14714
rect 1636 14662 1666 14714
rect 1666 14662 1678 14714
rect 1678 14662 1692 14714
rect 1716 14662 1730 14714
rect 1730 14662 1742 14714
rect 1742 14662 1772 14714
rect 1796 14662 1806 14714
rect 1806 14662 1852 14714
rect 1556 14660 1612 14662
rect 1636 14660 1692 14662
rect 1716 14660 1772 14662
rect 1796 14660 1852 14662
rect 5556 14714 5612 14716
rect 5636 14714 5692 14716
rect 5716 14714 5772 14716
rect 5796 14714 5852 14716
rect 5556 14662 5602 14714
rect 5602 14662 5612 14714
rect 5636 14662 5666 14714
rect 5666 14662 5678 14714
rect 5678 14662 5692 14714
rect 5716 14662 5730 14714
rect 5730 14662 5742 14714
rect 5742 14662 5772 14714
rect 5796 14662 5806 14714
rect 5806 14662 5852 14714
rect 5556 14660 5612 14662
rect 5636 14660 5692 14662
rect 5716 14660 5772 14662
rect 5796 14660 5852 14662
rect 9556 14714 9612 14716
rect 9636 14714 9692 14716
rect 9716 14714 9772 14716
rect 9796 14714 9852 14716
rect 9556 14662 9602 14714
rect 9602 14662 9612 14714
rect 9636 14662 9666 14714
rect 9666 14662 9678 14714
rect 9678 14662 9692 14714
rect 9716 14662 9730 14714
rect 9730 14662 9742 14714
rect 9742 14662 9772 14714
rect 9796 14662 9806 14714
rect 9806 14662 9852 14714
rect 9556 14660 9612 14662
rect 9636 14660 9692 14662
rect 9716 14660 9772 14662
rect 9796 14660 9852 14662
rect 13556 14714 13612 14716
rect 13636 14714 13692 14716
rect 13716 14714 13772 14716
rect 13796 14714 13852 14716
rect 13556 14662 13602 14714
rect 13602 14662 13612 14714
rect 13636 14662 13666 14714
rect 13666 14662 13678 14714
rect 13678 14662 13692 14714
rect 13716 14662 13730 14714
rect 13730 14662 13742 14714
rect 13742 14662 13772 14714
rect 13796 14662 13806 14714
rect 13806 14662 13852 14714
rect 13556 14660 13612 14662
rect 13636 14660 13692 14662
rect 13716 14660 13772 14662
rect 13796 14660 13852 14662
rect 17556 14714 17612 14716
rect 17636 14714 17692 14716
rect 17716 14714 17772 14716
rect 17796 14714 17852 14716
rect 17556 14662 17602 14714
rect 17602 14662 17612 14714
rect 17636 14662 17666 14714
rect 17666 14662 17678 14714
rect 17678 14662 17692 14714
rect 17716 14662 17730 14714
rect 17730 14662 17742 14714
rect 17742 14662 17772 14714
rect 17796 14662 17806 14714
rect 17806 14662 17852 14714
rect 17556 14660 17612 14662
rect 17636 14660 17692 14662
rect 17716 14660 17772 14662
rect 17796 14660 17852 14662
rect 2216 14170 2272 14172
rect 2296 14170 2352 14172
rect 2376 14170 2432 14172
rect 2456 14170 2512 14172
rect 2216 14118 2262 14170
rect 2262 14118 2272 14170
rect 2296 14118 2326 14170
rect 2326 14118 2338 14170
rect 2338 14118 2352 14170
rect 2376 14118 2390 14170
rect 2390 14118 2402 14170
rect 2402 14118 2432 14170
rect 2456 14118 2466 14170
rect 2466 14118 2512 14170
rect 2216 14116 2272 14118
rect 2296 14116 2352 14118
rect 2376 14116 2432 14118
rect 2456 14116 2512 14118
rect 6216 14170 6272 14172
rect 6296 14170 6352 14172
rect 6376 14170 6432 14172
rect 6456 14170 6512 14172
rect 6216 14118 6262 14170
rect 6262 14118 6272 14170
rect 6296 14118 6326 14170
rect 6326 14118 6338 14170
rect 6338 14118 6352 14170
rect 6376 14118 6390 14170
rect 6390 14118 6402 14170
rect 6402 14118 6432 14170
rect 6456 14118 6466 14170
rect 6466 14118 6512 14170
rect 6216 14116 6272 14118
rect 6296 14116 6352 14118
rect 6376 14116 6432 14118
rect 6456 14116 6512 14118
rect 10216 14170 10272 14172
rect 10296 14170 10352 14172
rect 10376 14170 10432 14172
rect 10456 14170 10512 14172
rect 10216 14118 10262 14170
rect 10262 14118 10272 14170
rect 10296 14118 10326 14170
rect 10326 14118 10338 14170
rect 10338 14118 10352 14170
rect 10376 14118 10390 14170
rect 10390 14118 10402 14170
rect 10402 14118 10432 14170
rect 10456 14118 10466 14170
rect 10466 14118 10512 14170
rect 10216 14116 10272 14118
rect 10296 14116 10352 14118
rect 10376 14116 10432 14118
rect 10456 14116 10512 14118
rect 14216 14170 14272 14172
rect 14296 14170 14352 14172
rect 14376 14170 14432 14172
rect 14456 14170 14512 14172
rect 14216 14118 14262 14170
rect 14262 14118 14272 14170
rect 14296 14118 14326 14170
rect 14326 14118 14338 14170
rect 14338 14118 14352 14170
rect 14376 14118 14390 14170
rect 14390 14118 14402 14170
rect 14402 14118 14432 14170
rect 14456 14118 14466 14170
rect 14466 14118 14512 14170
rect 14216 14116 14272 14118
rect 14296 14116 14352 14118
rect 14376 14116 14432 14118
rect 14456 14116 14512 14118
rect 18216 14170 18272 14172
rect 18296 14170 18352 14172
rect 18376 14170 18432 14172
rect 18456 14170 18512 14172
rect 18216 14118 18262 14170
rect 18262 14118 18272 14170
rect 18296 14118 18326 14170
rect 18326 14118 18338 14170
rect 18338 14118 18352 14170
rect 18376 14118 18390 14170
rect 18390 14118 18402 14170
rect 18402 14118 18432 14170
rect 18456 14118 18466 14170
rect 18466 14118 18512 14170
rect 18216 14116 18272 14118
rect 18296 14116 18352 14118
rect 18376 14116 18432 14118
rect 18456 14116 18512 14118
rect 1556 13626 1612 13628
rect 1636 13626 1692 13628
rect 1716 13626 1772 13628
rect 1796 13626 1852 13628
rect 1556 13574 1602 13626
rect 1602 13574 1612 13626
rect 1636 13574 1666 13626
rect 1666 13574 1678 13626
rect 1678 13574 1692 13626
rect 1716 13574 1730 13626
rect 1730 13574 1742 13626
rect 1742 13574 1772 13626
rect 1796 13574 1806 13626
rect 1806 13574 1852 13626
rect 1556 13572 1612 13574
rect 1636 13572 1692 13574
rect 1716 13572 1772 13574
rect 1796 13572 1852 13574
rect 5556 13626 5612 13628
rect 5636 13626 5692 13628
rect 5716 13626 5772 13628
rect 5796 13626 5852 13628
rect 5556 13574 5602 13626
rect 5602 13574 5612 13626
rect 5636 13574 5666 13626
rect 5666 13574 5678 13626
rect 5678 13574 5692 13626
rect 5716 13574 5730 13626
rect 5730 13574 5742 13626
rect 5742 13574 5772 13626
rect 5796 13574 5806 13626
rect 5806 13574 5852 13626
rect 5556 13572 5612 13574
rect 5636 13572 5692 13574
rect 5716 13572 5772 13574
rect 5796 13572 5852 13574
rect 9556 13626 9612 13628
rect 9636 13626 9692 13628
rect 9716 13626 9772 13628
rect 9796 13626 9852 13628
rect 9556 13574 9602 13626
rect 9602 13574 9612 13626
rect 9636 13574 9666 13626
rect 9666 13574 9678 13626
rect 9678 13574 9692 13626
rect 9716 13574 9730 13626
rect 9730 13574 9742 13626
rect 9742 13574 9772 13626
rect 9796 13574 9806 13626
rect 9806 13574 9852 13626
rect 9556 13572 9612 13574
rect 9636 13572 9692 13574
rect 9716 13572 9772 13574
rect 9796 13572 9852 13574
rect 13556 13626 13612 13628
rect 13636 13626 13692 13628
rect 13716 13626 13772 13628
rect 13796 13626 13852 13628
rect 13556 13574 13602 13626
rect 13602 13574 13612 13626
rect 13636 13574 13666 13626
rect 13666 13574 13678 13626
rect 13678 13574 13692 13626
rect 13716 13574 13730 13626
rect 13730 13574 13742 13626
rect 13742 13574 13772 13626
rect 13796 13574 13806 13626
rect 13806 13574 13852 13626
rect 13556 13572 13612 13574
rect 13636 13572 13692 13574
rect 13716 13572 13772 13574
rect 13796 13572 13852 13574
rect 17556 13626 17612 13628
rect 17636 13626 17692 13628
rect 17716 13626 17772 13628
rect 17796 13626 17852 13628
rect 17556 13574 17602 13626
rect 17602 13574 17612 13626
rect 17636 13574 17666 13626
rect 17666 13574 17678 13626
rect 17678 13574 17692 13626
rect 17716 13574 17730 13626
rect 17730 13574 17742 13626
rect 17742 13574 17772 13626
rect 17796 13574 17806 13626
rect 17806 13574 17852 13626
rect 17556 13572 17612 13574
rect 17636 13572 17692 13574
rect 17716 13572 17772 13574
rect 17796 13572 17852 13574
rect 2216 13082 2272 13084
rect 2296 13082 2352 13084
rect 2376 13082 2432 13084
rect 2456 13082 2512 13084
rect 2216 13030 2262 13082
rect 2262 13030 2272 13082
rect 2296 13030 2326 13082
rect 2326 13030 2338 13082
rect 2338 13030 2352 13082
rect 2376 13030 2390 13082
rect 2390 13030 2402 13082
rect 2402 13030 2432 13082
rect 2456 13030 2466 13082
rect 2466 13030 2512 13082
rect 2216 13028 2272 13030
rect 2296 13028 2352 13030
rect 2376 13028 2432 13030
rect 2456 13028 2512 13030
rect 6216 13082 6272 13084
rect 6296 13082 6352 13084
rect 6376 13082 6432 13084
rect 6456 13082 6512 13084
rect 6216 13030 6262 13082
rect 6262 13030 6272 13082
rect 6296 13030 6326 13082
rect 6326 13030 6338 13082
rect 6338 13030 6352 13082
rect 6376 13030 6390 13082
rect 6390 13030 6402 13082
rect 6402 13030 6432 13082
rect 6456 13030 6466 13082
rect 6466 13030 6512 13082
rect 6216 13028 6272 13030
rect 6296 13028 6352 13030
rect 6376 13028 6432 13030
rect 6456 13028 6512 13030
rect 10216 13082 10272 13084
rect 10296 13082 10352 13084
rect 10376 13082 10432 13084
rect 10456 13082 10512 13084
rect 10216 13030 10262 13082
rect 10262 13030 10272 13082
rect 10296 13030 10326 13082
rect 10326 13030 10338 13082
rect 10338 13030 10352 13082
rect 10376 13030 10390 13082
rect 10390 13030 10402 13082
rect 10402 13030 10432 13082
rect 10456 13030 10466 13082
rect 10466 13030 10512 13082
rect 10216 13028 10272 13030
rect 10296 13028 10352 13030
rect 10376 13028 10432 13030
rect 10456 13028 10512 13030
rect 14216 13082 14272 13084
rect 14296 13082 14352 13084
rect 14376 13082 14432 13084
rect 14456 13082 14512 13084
rect 14216 13030 14262 13082
rect 14262 13030 14272 13082
rect 14296 13030 14326 13082
rect 14326 13030 14338 13082
rect 14338 13030 14352 13082
rect 14376 13030 14390 13082
rect 14390 13030 14402 13082
rect 14402 13030 14432 13082
rect 14456 13030 14466 13082
rect 14466 13030 14512 13082
rect 14216 13028 14272 13030
rect 14296 13028 14352 13030
rect 14376 13028 14432 13030
rect 14456 13028 14512 13030
rect 18216 13082 18272 13084
rect 18296 13082 18352 13084
rect 18376 13082 18432 13084
rect 18456 13082 18512 13084
rect 18216 13030 18262 13082
rect 18262 13030 18272 13082
rect 18296 13030 18326 13082
rect 18326 13030 18338 13082
rect 18338 13030 18352 13082
rect 18376 13030 18390 13082
rect 18390 13030 18402 13082
rect 18402 13030 18432 13082
rect 18456 13030 18466 13082
rect 18466 13030 18512 13082
rect 18216 13028 18272 13030
rect 18296 13028 18352 13030
rect 18376 13028 18432 13030
rect 18456 13028 18512 13030
rect 1556 12538 1612 12540
rect 1636 12538 1692 12540
rect 1716 12538 1772 12540
rect 1796 12538 1852 12540
rect 1556 12486 1602 12538
rect 1602 12486 1612 12538
rect 1636 12486 1666 12538
rect 1666 12486 1678 12538
rect 1678 12486 1692 12538
rect 1716 12486 1730 12538
rect 1730 12486 1742 12538
rect 1742 12486 1772 12538
rect 1796 12486 1806 12538
rect 1806 12486 1852 12538
rect 1556 12484 1612 12486
rect 1636 12484 1692 12486
rect 1716 12484 1772 12486
rect 1796 12484 1852 12486
rect 5556 12538 5612 12540
rect 5636 12538 5692 12540
rect 5716 12538 5772 12540
rect 5796 12538 5852 12540
rect 5556 12486 5602 12538
rect 5602 12486 5612 12538
rect 5636 12486 5666 12538
rect 5666 12486 5678 12538
rect 5678 12486 5692 12538
rect 5716 12486 5730 12538
rect 5730 12486 5742 12538
rect 5742 12486 5772 12538
rect 5796 12486 5806 12538
rect 5806 12486 5852 12538
rect 5556 12484 5612 12486
rect 5636 12484 5692 12486
rect 5716 12484 5772 12486
rect 5796 12484 5852 12486
rect 9556 12538 9612 12540
rect 9636 12538 9692 12540
rect 9716 12538 9772 12540
rect 9796 12538 9852 12540
rect 9556 12486 9602 12538
rect 9602 12486 9612 12538
rect 9636 12486 9666 12538
rect 9666 12486 9678 12538
rect 9678 12486 9692 12538
rect 9716 12486 9730 12538
rect 9730 12486 9742 12538
rect 9742 12486 9772 12538
rect 9796 12486 9806 12538
rect 9806 12486 9852 12538
rect 9556 12484 9612 12486
rect 9636 12484 9692 12486
rect 9716 12484 9772 12486
rect 9796 12484 9852 12486
rect 13556 12538 13612 12540
rect 13636 12538 13692 12540
rect 13716 12538 13772 12540
rect 13796 12538 13852 12540
rect 13556 12486 13602 12538
rect 13602 12486 13612 12538
rect 13636 12486 13666 12538
rect 13666 12486 13678 12538
rect 13678 12486 13692 12538
rect 13716 12486 13730 12538
rect 13730 12486 13742 12538
rect 13742 12486 13772 12538
rect 13796 12486 13806 12538
rect 13806 12486 13852 12538
rect 13556 12484 13612 12486
rect 13636 12484 13692 12486
rect 13716 12484 13772 12486
rect 13796 12484 13852 12486
rect 17556 12538 17612 12540
rect 17636 12538 17692 12540
rect 17716 12538 17772 12540
rect 17796 12538 17852 12540
rect 17556 12486 17602 12538
rect 17602 12486 17612 12538
rect 17636 12486 17666 12538
rect 17666 12486 17678 12538
rect 17678 12486 17692 12538
rect 17716 12486 17730 12538
rect 17730 12486 17742 12538
rect 17742 12486 17772 12538
rect 17796 12486 17806 12538
rect 17806 12486 17852 12538
rect 17556 12484 17612 12486
rect 17636 12484 17692 12486
rect 17716 12484 17772 12486
rect 17796 12484 17852 12486
rect 2216 11994 2272 11996
rect 2296 11994 2352 11996
rect 2376 11994 2432 11996
rect 2456 11994 2512 11996
rect 2216 11942 2262 11994
rect 2262 11942 2272 11994
rect 2296 11942 2326 11994
rect 2326 11942 2338 11994
rect 2338 11942 2352 11994
rect 2376 11942 2390 11994
rect 2390 11942 2402 11994
rect 2402 11942 2432 11994
rect 2456 11942 2466 11994
rect 2466 11942 2512 11994
rect 2216 11940 2272 11942
rect 2296 11940 2352 11942
rect 2376 11940 2432 11942
rect 2456 11940 2512 11942
rect 6216 11994 6272 11996
rect 6296 11994 6352 11996
rect 6376 11994 6432 11996
rect 6456 11994 6512 11996
rect 6216 11942 6262 11994
rect 6262 11942 6272 11994
rect 6296 11942 6326 11994
rect 6326 11942 6338 11994
rect 6338 11942 6352 11994
rect 6376 11942 6390 11994
rect 6390 11942 6402 11994
rect 6402 11942 6432 11994
rect 6456 11942 6466 11994
rect 6466 11942 6512 11994
rect 6216 11940 6272 11942
rect 6296 11940 6352 11942
rect 6376 11940 6432 11942
rect 6456 11940 6512 11942
rect 10216 11994 10272 11996
rect 10296 11994 10352 11996
rect 10376 11994 10432 11996
rect 10456 11994 10512 11996
rect 10216 11942 10262 11994
rect 10262 11942 10272 11994
rect 10296 11942 10326 11994
rect 10326 11942 10338 11994
rect 10338 11942 10352 11994
rect 10376 11942 10390 11994
rect 10390 11942 10402 11994
rect 10402 11942 10432 11994
rect 10456 11942 10466 11994
rect 10466 11942 10512 11994
rect 10216 11940 10272 11942
rect 10296 11940 10352 11942
rect 10376 11940 10432 11942
rect 10456 11940 10512 11942
rect 14216 11994 14272 11996
rect 14296 11994 14352 11996
rect 14376 11994 14432 11996
rect 14456 11994 14512 11996
rect 14216 11942 14262 11994
rect 14262 11942 14272 11994
rect 14296 11942 14326 11994
rect 14326 11942 14338 11994
rect 14338 11942 14352 11994
rect 14376 11942 14390 11994
rect 14390 11942 14402 11994
rect 14402 11942 14432 11994
rect 14456 11942 14466 11994
rect 14466 11942 14512 11994
rect 14216 11940 14272 11942
rect 14296 11940 14352 11942
rect 14376 11940 14432 11942
rect 14456 11940 14512 11942
rect 18216 11994 18272 11996
rect 18296 11994 18352 11996
rect 18376 11994 18432 11996
rect 18456 11994 18512 11996
rect 18216 11942 18262 11994
rect 18262 11942 18272 11994
rect 18296 11942 18326 11994
rect 18326 11942 18338 11994
rect 18338 11942 18352 11994
rect 18376 11942 18390 11994
rect 18390 11942 18402 11994
rect 18402 11942 18432 11994
rect 18456 11942 18466 11994
rect 18466 11942 18512 11994
rect 18216 11940 18272 11942
rect 18296 11940 18352 11942
rect 18376 11940 18432 11942
rect 18456 11940 18512 11942
rect 846 11772 848 11792
rect 848 11772 900 11792
rect 900 11772 902 11792
rect 846 11736 902 11772
rect 1556 11450 1612 11452
rect 1636 11450 1692 11452
rect 1716 11450 1772 11452
rect 1796 11450 1852 11452
rect 1556 11398 1602 11450
rect 1602 11398 1612 11450
rect 1636 11398 1666 11450
rect 1666 11398 1678 11450
rect 1678 11398 1692 11450
rect 1716 11398 1730 11450
rect 1730 11398 1742 11450
rect 1742 11398 1772 11450
rect 1796 11398 1806 11450
rect 1806 11398 1852 11450
rect 1556 11396 1612 11398
rect 1636 11396 1692 11398
rect 1716 11396 1772 11398
rect 1796 11396 1852 11398
rect 5556 11450 5612 11452
rect 5636 11450 5692 11452
rect 5716 11450 5772 11452
rect 5796 11450 5852 11452
rect 5556 11398 5602 11450
rect 5602 11398 5612 11450
rect 5636 11398 5666 11450
rect 5666 11398 5678 11450
rect 5678 11398 5692 11450
rect 5716 11398 5730 11450
rect 5730 11398 5742 11450
rect 5742 11398 5772 11450
rect 5796 11398 5806 11450
rect 5806 11398 5852 11450
rect 5556 11396 5612 11398
rect 5636 11396 5692 11398
rect 5716 11396 5772 11398
rect 5796 11396 5852 11398
rect 9556 11450 9612 11452
rect 9636 11450 9692 11452
rect 9716 11450 9772 11452
rect 9796 11450 9852 11452
rect 9556 11398 9602 11450
rect 9602 11398 9612 11450
rect 9636 11398 9666 11450
rect 9666 11398 9678 11450
rect 9678 11398 9692 11450
rect 9716 11398 9730 11450
rect 9730 11398 9742 11450
rect 9742 11398 9772 11450
rect 9796 11398 9806 11450
rect 9806 11398 9852 11450
rect 9556 11396 9612 11398
rect 9636 11396 9692 11398
rect 9716 11396 9772 11398
rect 9796 11396 9852 11398
rect 13556 11450 13612 11452
rect 13636 11450 13692 11452
rect 13716 11450 13772 11452
rect 13796 11450 13852 11452
rect 13556 11398 13602 11450
rect 13602 11398 13612 11450
rect 13636 11398 13666 11450
rect 13666 11398 13678 11450
rect 13678 11398 13692 11450
rect 13716 11398 13730 11450
rect 13730 11398 13742 11450
rect 13742 11398 13772 11450
rect 13796 11398 13806 11450
rect 13806 11398 13852 11450
rect 13556 11396 13612 11398
rect 13636 11396 13692 11398
rect 13716 11396 13772 11398
rect 13796 11396 13852 11398
rect 17556 11450 17612 11452
rect 17636 11450 17692 11452
rect 17716 11450 17772 11452
rect 17796 11450 17852 11452
rect 17556 11398 17602 11450
rect 17602 11398 17612 11450
rect 17636 11398 17666 11450
rect 17666 11398 17678 11450
rect 17678 11398 17692 11450
rect 17716 11398 17730 11450
rect 17730 11398 17742 11450
rect 17742 11398 17772 11450
rect 17796 11398 17806 11450
rect 17806 11398 17852 11450
rect 17556 11396 17612 11398
rect 17636 11396 17692 11398
rect 17716 11396 17772 11398
rect 17796 11396 17852 11398
rect 1398 10920 1454 10976
rect 2216 10906 2272 10908
rect 2296 10906 2352 10908
rect 2376 10906 2432 10908
rect 2456 10906 2512 10908
rect 2216 10854 2262 10906
rect 2262 10854 2272 10906
rect 2296 10854 2326 10906
rect 2326 10854 2338 10906
rect 2338 10854 2352 10906
rect 2376 10854 2390 10906
rect 2390 10854 2402 10906
rect 2402 10854 2432 10906
rect 2456 10854 2466 10906
rect 2466 10854 2512 10906
rect 2216 10852 2272 10854
rect 2296 10852 2352 10854
rect 2376 10852 2432 10854
rect 2456 10852 2512 10854
rect 6216 10906 6272 10908
rect 6296 10906 6352 10908
rect 6376 10906 6432 10908
rect 6456 10906 6512 10908
rect 6216 10854 6262 10906
rect 6262 10854 6272 10906
rect 6296 10854 6326 10906
rect 6326 10854 6338 10906
rect 6338 10854 6352 10906
rect 6376 10854 6390 10906
rect 6390 10854 6402 10906
rect 6402 10854 6432 10906
rect 6456 10854 6466 10906
rect 6466 10854 6512 10906
rect 6216 10852 6272 10854
rect 6296 10852 6352 10854
rect 6376 10852 6432 10854
rect 6456 10852 6512 10854
rect 10216 10906 10272 10908
rect 10296 10906 10352 10908
rect 10376 10906 10432 10908
rect 10456 10906 10512 10908
rect 10216 10854 10262 10906
rect 10262 10854 10272 10906
rect 10296 10854 10326 10906
rect 10326 10854 10338 10906
rect 10338 10854 10352 10906
rect 10376 10854 10390 10906
rect 10390 10854 10402 10906
rect 10402 10854 10432 10906
rect 10456 10854 10466 10906
rect 10466 10854 10512 10906
rect 10216 10852 10272 10854
rect 10296 10852 10352 10854
rect 10376 10852 10432 10854
rect 10456 10852 10512 10854
rect 14216 10906 14272 10908
rect 14296 10906 14352 10908
rect 14376 10906 14432 10908
rect 14456 10906 14512 10908
rect 14216 10854 14262 10906
rect 14262 10854 14272 10906
rect 14296 10854 14326 10906
rect 14326 10854 14338 10906
rect 14338 10854 14352 10906
rect 14376 10854 14390 10906
rect 14390 10854 14402 10906
rect 14402 10854 14432 10906
rect 14456 10854 14466 10906
rect 14466 10854 14512 10906
rect 14216 10852 14272 10854
rect 14296 10852 14352 10854
rect 14376 10852 14432 10854
rect 14456 10852 14512 10854
rect 18216 10906 18272 10908
rect 18296 10906 18352 10908
rect 18376 10906 18432 10908
rect 18456 10906 18512 10908
rect 18216 10854 18262 10906
rect 18262 10854 18272 10906
rect 18296 10854 18326 10906
rect 18326 10854 18338 10906
rect 18338 10854 18352 10906
rect 18376 10854 18390 10906
rect 18390 10854 18402 10906
rect 18402 10854 18432 10906
rect 18456 10854 18466 10906
rect 18466 10854 18512 10906
rect 18216 10852 18272 10854
rect 18296 10852 18352 10854
rect 18376 10852 18432 10854
rect 18456 10852 18512 10854
rect 846 10412 848 10432
rect 848 10412 900 10432
rect 900 10412 902 10432
rect 846 10376 902 10412
rect 1556 10362 1612 10364
rect 1636 10362 1692 10364
rect 1716 10362 1772 10364
rect 1796 10362 1852 10364
rect 1556 10310 1602 10362
rect 1602 10310 1612 10362
rect 1636 10310 1666 10362
rect 1666 10310 1678 10362
rect 1678 10310 1692 10362
rect 1716 10310 1730 10362
rect 1730 10310 1742 10362
rect 1742 10310 1772 10362
rect 1796 10310 1806 10362
rect 1806 10310 1852 10362
rect 1556 10308 1612 10310
rect 1636 10308 1692 10310
rect 1716 10308 1772 10310
rect 1796 10308 1852 10310
rect 5556 10362 5612 10364
rect 5636 10362 5692 10364
rect 5716 10362 5772 10364
rect 5796 10362 5852 10364
rect 5556 10310 5602 10362
rect 5602 10310 5612 10362
rect 5636 10310 5666 10362
rect 5666 10310 5678 10362
rect 5678 10310 5692 10362
rect 5716 10310 5730 10362
rect 5730 10310 5742 10362
rect 5742 10310 5772 10362
rect 5796 10310 5806 10362
rect 5806 10310 5852 10362
rect 5556 10308 5612 10310
rect 5636 10308 5692 10310
rect 5716 10308 5772 10310
rect 5796 10308 5852 10310
rect 9556 10362 9612 10364
rect 9636 10362 9692 10364
rect 9716 10362 9772 10364
rect 9796 10362 9852 10364
rect 9556 10310 9602 10362
rect 9602 10310 9612 10362
rect 9636 10310 9666 10362
rect 9666 10310 9678 10362
rect 9678 10310 9692 10362
rect 9716 10310 9730 10362
rect 9730 10310 9742 10362
rect 9742 10310 9772 10362
rect 9796 10310 9806 10362
rect 9806 10310 9852 10362
rect 9556 10308 9612 10310
rect 9636 10308 9692 10310
rect 9716 10308 9772 10310
rect 9796 10308 9852 10310
rect 13556 10362 13612 10364
rect 13636 10362 13692 10364
rect 13716 10362 13772 10364
rect 13796 10362 13852 10364
rect 13556 10310 13602 10362
rect 13602 10310 13612 10362
rect 13636 10310 13666 10362
rect 13666 10310 13678 10362
rect 13678 10310 13692 10362
rect 13716 10310 13730 10362
rect 13730 10310 13742 10362
rect 13742 10310 13772 10362
rect 13796 10310 13806 10362
rect 13806 10310 13852 10362
rect 13556 10308 13612 10310
rect 13636 10308 13692 10310
rect 13716 10308 13772 10310
rect 13796 10308 13852 10310
rect 17556 10362 17612 10364
rect 17636 10362 17692 10364
rect 17716 10362 17772 10364
rect 17796 10362 17852 10364
rect 17556 10310 17602 10362
rect 17602 10310 17612 10362
rect 17636 10310 17666 10362
rect 17666 10310 17678 10362
rect 17678 10310 17692 10362
rect 17716 10310 17730 10362
rect 17730 10310 17742 10362
rect 17742 10310 17772 10362
rect 17796 10310 17806 10362
rect 17806 10310 17852 10362
rect 17556 10308 17612 10310
rect 17636 10308 17692 10310
rect 17716 10308 17772 10310
rect 17796 10308 17852 10310
rect 18510 10240 18566 10296
rect 2216 9818 2272 9820
rect 2296 9818 2352 9820
rect 2376 9818 2432 9820
rect 2456 9818 2512 9820
rect 2216 9766 2262 9818
rect 2262 9766 2272 9818
rect 2296 9766 2326 9818
rect 2326 9766 2338 9818
rect 2338 9766 2352 9818
rect 2376 9766 2390 9818
rect 2390 9766 2402 9818
rect 2402 9766 2432 9818
rect 2456 9766 2466 9818
rect 2466 9766 2512 9818
rect 2216 9764 2272 9766
rect 2296 9764 2352 9766
rect 2376 9764 2432 9766
rect 2456 9764 2512 9766
rect 6216 9818 6272 9820
rect 6296 9818 6352 9820
rect 6376 9818 6432 9820
rect 6456 9818 6512 9820
rect 6216 9766 6262 9818
rect 6262 9766 6272 9818
rect 6296 9766 6326 9818
rect 6326 9766 6338 9818
rect 6338 9766 6352 9818
rect 6376 9766 6390 9818
rect 6390 9766 6402 9818
rect 6402 9766 6432 9818
rect 6456 9766 6466 9818
rect 6466 9766 6512 9818
rect 6216 9764 6272 9766
rect 6296 9764 6352 9766
rect 6376 9764 6432 9766
rect 6456 9764 6512 9766
rect 10216 9818 10272 9820
rect 10296 9818 10352 9820
rect 10376 9818 10432 9820
rect 10456 9818 10512 9820
rect 10216 9766 10262 9818
rect 10262 9766 10272 9818
rect 10296 9766 10326 9818
rect 10326 9766 10338 9818
rect 10338 9766 10352 9818
rect 10376 9766 10390 9818
rect 10390 9766 10402 9818
rect 10402 9766 10432 9818
rect 10456 9766 10466 9818
rect 10466 9766 10512 9818
rect 10216 9764 10272 9766
rect 10296 9764 10352 9766
rect 10376 9764 10432 9766
rect 10456 9764 10512 9766
rect 14216 9818 14272 9820
rect 14296 9818 14352 9820
rect 14376 9818 14432 9820
rect 14456 9818 14512 9820
rect 14216 9766 14262 9818
rect 14262 9766 14272 9818
rect 14296 9766 14326 9818
rect 14326 9766 14338 9818
rect 14338 9766 14352 9818
rect 14376 9766 14390 9818
rect 14390 9766 14402 9818
rect 14402 9766 14432 9818
rect 14456 9766 14466 9818
rect 14466 9766 14512 9818
rect 14216 9764 14272 9766
rect 14296 9764 14352 9766
rect 14376 9764 14432 9766
rect 14456 9764 14512 9766
rect 18216 9818 18272 9820
rect 18296 9818 18352 9820
rect 18376 9818 18432 9820
rect 18456 9818 18512 9820
rect 18216 9766 18262 9818
rect 18262 9766 18272 9818
rect 18296 9766 18326 9818
rect 18326 9766 18338 9818
rect 18338 9766 18352 9818
rect 18376 9766 18390 9818
rect 18390 9766 18402 9818
rect 18402 9766 18432 9818
rect 18456 9766 18466 9818
rect 18466 9766 18512 9818
rect 18216 9764 18272 9766
rect 18296 9764 18352 9766
rect 18376 9764 18432 9766
rect 18456 9764 18512 9766
rect 1398 9560 1454 9616
rect 1556 9274 1612 9276
rect 1636 9274 1692 9276
rect 1716 9274 1772 9276
rect 1796 9274 1852 9276
rect 1556 9222 1602 9274
rect 1602 9222 1612 9274
rect 1636 9222 1666 9274
rect 1666 9222 1678 9274
rect 1678 9222 1692 9274
rect 1716 9222 1730 9274
rect 1730 9222 1742 9274
rect 1742 9222 1772 9274
rect 1796 9222 1806 9274
rect 1806 9222 1852 9274
rect 1556 9220 1612 9222
rect 1636 9220 1692 9222
rect 1716 9220 1772 9222
rect 1796 9220 1852 9222
rect 5556 9274 5612 9276
rect 5636 9274 5692 9276
rect 5716 9274 5772 9276
rect 5796 9274 5852 9276
rect 5556 9222 5602 9274
rect 5602 9222 5612 9274
rect 5636 9222 5666 9274
rect 5666 9222 5678 9274
rect 5678 9222 5692 9274
rect 5716 9222 5730 9274
rect 5730 9222 5742 9274
rect 5742 9222 5772 9274
rect 5796 9222 5806 9274
rect 5806 9222 5852 9274
rect 5556 9220 5612 9222
rect 5636 9220 5692 9222
rect 5716 9220 5772 9222
rect 5796 9220 5852 9222
rect 9556 9274 9612 9276
rect 9636 9274 9692 9276
rect 9716 9274 9772 9276
rect 9796 9274 9852 9276
rect 9556 9222 9602 9274
rect 9602 9222 9612 9274
rect 9636 9222 9666 9274
rect 9666 9222 9678 9274
rect 9678 9222 9692 9274
rect 9716 9222 9730 9274
rect 9730 9222 9742 9274
rect 9742 9222 9772 9274
rect 9796 9222 9806 9274
rect 9806 9222 9852 9274
rect 9556 9220 9612 9222
rect 9636 9220 9692 9222
rect 9716 9220 9772 9222
rect 9796 9220 9852 9222
rect 13556 9274 13612 9276
rect 13636 9274 13692 9276
rect 13716 9274 13772 9276
rect 13796 9274 13852 9276
rect 13556 9222 13602 9274
rect 13602 9222 13612 9274
rect 13636 9222 13666 9274
rect 13666 9222 13678 9274
rect 13678 9222 13692 9274
rect 13716 9222 13730 9274
rect 13730 9222 13742 9274
rect 13742 9222 13772 9274
rect 13796 9222 13806 9274
rect 13806 9222 13852 9274
rect 13556 9220 13612 9222
rect 13636 9220 13692 9222
rect 13716 9220 13772 9222
rect 13796 9220 13852 9222
rect 17556 9274 17612 9276
rect 17636 9274 17692 9276
rect 17716 9274 17772 9276
rect 17796 9274 17852 9276
rect 17556 9222 17602 9274
rect 17602 9222 17612 9274
rect 17636 9222 17666 9274
rect 17666 9222 17678 9274
rect 17678 9222 17692 9274
rect 17716 9222 17730 9274
rect 17730 9222 17742 9274
rect 17742 9222 17772 9274
rect 17796 9222 17806 9274
rect 17806 9222 17852 9274
rect 17556 9220 17612 9222
rect 17636 9220 17692 9222
rect 17716 9220 17772 9222
rect 17796 9220 17852 9222
rect 846 9036 902 9072
rect 846 9016 848 9036
rect 848 9016 900 9036
rect 900 9016 902 9036
rect 2216 8730 2272 8732
rect 2296 8730 2352 8732
rect 2376 8730 2432 8732
rect 2456 8730 2512 8732
rect 2216 8678 2262 8730
rect 2262 8678 2272 8730
rect 2296 8678 2326 8730
rect 2326 8678 2338 8730
rect 2338 8678 2352 8730
rect 2376 8678 2390 8730
rect 2390 8678 2402 8730
rect 2402 8678 2432 8730
rect 2456 8678 2466 8730
rect 2466 8678 2512 8730
rect 2216 8676 2272 8678
rect 2296 8676 2352 8678
rect 2376 8676 2432 8678
rect 2456 8676 2512 8678
rect 6216 8730 6272 8732
rect 6296 8730 6352 8732
rect 6376 8730 6432 8732
rect 6456 8730 6512 8732
rect 6216 8678 6262 8730
rect 6262 8678 6272 8730
rect 6296 8678 6326 8730
rect 6326 8678 6338 8730
rect 6338 8678 6352 8730
rect 6376 8678 6390 8730
rect 6390 8678 6402 8730
rect 6402 8678 6432 8730
rect 6456 8678 6466 8730
rect 6466 8678 6512 8730
rect 6216 8676 6272 8678
rect 6296 8676 6352 8678
rect 6376 8676 6432 8678
rect 6456 8676 6512 8678
rect 10216 8730 10272 8732
rect 10296 8730 10352 8732
rect 10376 8730 10432 8732
rect 10456 8730 10512 8732
rect 10216 8678 10262 8730
rect 10262 8678 10272 8730
rect 10296 8678 10326 8730
rect 10326 8678 10338 8730
rect 10338 8678 10352 8730
rect 10376 8678 10390 8730
rect 10390 8678 10402 8730
rect 10402 8678 10432 8730
rect 10456 8678 10466 8730
rect 10466 8678 10512 8730
rect 10216 8676 10272 8678
rect 10296 8676 10352 8678
rect 10376 8676 10432 8678
rect 10456 8676 10512 8678
rect 14216 8730 14272 8732
rect 14296 8730 14352 8732
rect 14376 8730 14432 8732
rect 14456 8730 14512 8732
rect 14216 8678 14262 8730
rect 14262 8678 14272 8730
rect 14296 8678 14326 8730
rect 14326 8678 14338 8730
rect 14338 8678 14352 8730
rect 14376 8678 14390 8730
rect 14390 8678 14402 8730
rect 14402 8678 14432 8730
rect 14456 8678 14466 8730
rect 14466 8678 14512 8730
rect 14216 8676 14272 8678
rect 14296 8676 14352 8678
rect 14376 8676 14432 8678
rect 14456 8676 14512 8678
rect 18216 8730 18272 8732
rect 18296 8730 18352 8732
rect 18376 8730 18432 8732
rect 18456 8730 18512 8732
rect 18216 8678 18262 8730
rect 18262 8678 18272 8730
rect 18296 8678 18326 8730
rect 18326 8678 18338 8730
rect 18338 8678 18352 8730
rect 18376 8678 18390 8730
rect 18390 8678 18402 8730
rect 18402 8678 18432 8730
rect 18456 8678 18466 8730
rect 18466 8678 18512 8730
rect 18216 8676 18272 8678
rect 18296 8676 18352 8678
rect 18376 8676 18432 8678
rect 18456 8676 18512 8678
rect 1398 8200 1454 8256
rect 1556 8186 1612 8188
rect 1636 8186 1692 8188
rect 1716 8186 1772 8188
rect 1796 8186 1852 8188
rect 1556 8134 1602 8186
rect 1602 8134 1612 8186
rect 1636 8134 1666 8186
rect 1666 8134 1678 8186
rect 1678 8134 1692 8186
rect 1716 8134 1730 8186
rect 1730 8134 1742 8186
rect 1742 8134 1772 8186
rect 1796 8134 1806 8186
rect 1806 8134 1852 8186
rect 1556 8132 1612 8134
rect 1636 8132 1692 8134
rect 1716 8132 1772 8134
rect 1796 8132 1852 8134
rect 5556 8186 5612 8188
rect 5636 8186 5692 8188
rect 5716 8186 5772 8188
rect 5796 8186 5852 8188
rect 5556 8134 5602 8186
rect 5602 8134 5612 8186
rect 5636 8134 5666 8186
rect 5666 8134 5678 8186
rect 5678 8134 5692 8186
rect 5716 8134 5730 8186
rect 5730 8134 5742 8186
rect 5742 8134 5772 8186
rect 5796 8134 5806 8186
rect 5806 8134 5852 8186
rect 5556 8132 5612 8134
rect 5636 8132 5692 8134
rect 5716 8132 5772 8134
rect 5796 8132 5852 8134
rect 9556 8186 9612 8188
rect 9636 8186 9692 8188
rect 9716 8186 9772 8188
rect 9796 8186 9852 8188
rect 9556 8134 9602 8186
rect 9602 8134 9612 8186
rect 9636 8134 9666 8186
rect 9666 8134 9678 8186
rect 9678 8134 9692 8186
rect 9716 8134 9730 8186
rect 9730 8134 9742 8186
rect 9742 8134 9772 8186
rect 9796 8134 9806 8186
rect 9806 8134 9852 8186
rect 9556 8132 9612 8134
rect 9636 8132 9692 8134
rect 9716 8132 9772 8134
rect 9796 8132 9852 8134
rect 13556 8186 13612 8188
rect 13636 8186 13692 8188
rect 13716 8186 13772 8188
rect 13796 8186 13852 8188
rect 13556 8134 13602 8186
rect 13602 8134 13612 8186
rect 13636 8134 13666 8186
rect 13666 8134 13678 8186
rect 13678 8134 13692 8186
rect 13716 8134 13730 8186
rect 13730 8134 13742 8186
rect 13742 8134 13772 8186
rect 13796 8134 13806 8186
rect 13806 8134 13852 8186
rect 13556 8132 13612 8134
rect 13636 8132 13692 8134
rect 13716 8132 13772 8134
rect 13796 8132 13852 8134
rect 17556 8186 17612 8188
rect 17636 8186 17692 8188
rect 17716 8186 17772 8188
rect 17796 8186 17852 8188
rect 17556 8134 17602 8186
rect 17602 8134 17612 8186
rect 17636 8134 17666 8186
rect 17666 8134 17678 8186
rect 17678 8134 17692 8186
rect 17716 8134 17730 8186
rect 17730 8134 17742 8186
rect 17742 8134 17772 8186
rect 17796 8134 17806 8186
rect 17806 8134 17852 8186
rect 17556 8132 17612 8134
rect 17636 8132 17692 8134
rect 17716 8132 17772 8134
rect 17796 8132 17852 8134
rect 2216 7642 2272 7644
rect 2296 7642 2352 7644
rect 2376 7642 2432 7644
rect 2456 7642 2512 7644
rect 2216 7590 2262 7642
rect 2262 7590 2272 7642
rect 2296 7590 2326 7642
rect 2326 7590 2338 7642
rect 2338 7590 2352 7642
rect 2376 7590 2390 7642
rect 2390 7590 2402 7642
rect 2402 7590 2432 7642
rect 2456 7590 2466 7642
rect 2466 7590 2512 7642
rect 2216 7588 2272 7590
rect 2296 7588 2352 7590
rect 2376 7588 2432 7590
rect 2456 7588 2512 7590
rect 6216 7642 6272 7644
rect 6296 7642 6352 7644
rect 6376 7642 6432 7644
rect 6456 7642 6512 7644
rect 6216 7590 6262 7642
rect 6262 7590 6272 7642
rect 6296 7590 6326 7642
rect 6326 7590 6338 7642
rect 6338 7590 6352 7642
rect 6376 7590 6390 7642
rect 6390 7590 6402 7642
rect 6402 7590 6432 7642
rect 6456 7590 6466 7642
rect 6466 7590 6512 7642
rect 6216 7588 6272 7590
rect 6296 7588 6352 7590
rect 6376 7588 6432 7590
rect 6456 7588 6512 7590
rect 10216 7642 10272 7644
rect 10296 7642 10352 7644
rect 10376 7642 10432 7644
rect 10456 7642 10512 7644
rect 10216 7590 10262 7642
rect 10262 7590 10272 7642
rect 10296 7590 10326 7642
rect 10326 7590 10338 7642
rect 10338 7590 10352 7642
rect 10376 7590 10390 7642
rect 10390 7590 10402 7642
rect 10402 7590 10432 7642
rect 10456 7590 10466 7642
rect 10466 7590 10512 7642
rect 10216 7588 10272 7590
rect 10296 7588 10352 7590
rect 10376 7588 10432 7590
rect 10456 7588 10512 7590
rect 14216 7642 14272 7644
rect 14296 7642 14352 7644
rect 14376 7642 14432 7644
rect 14456 7642 14512 7644
rect 14216 7590 14262 7642
rect 14262 7590 14272 7642
rect 14296 7590 14326 7642
rect 14326 7590 14338 7642
rect 14338 7590 14352 7642
rect 14376 7590 14390 7642
rect 14390 7590 14402 7642
rect 14402 7590 14432 7642
rect 14456 7590 14466 7642
rect 14466 7590 14512 7642
rect 14216 7588 14272 7590
rect 14296 7588 14352 7590
rect 14376 7588 14432 7590
rect 14456 7588 14512 7590
rect 18216 7642 18272 7644
rect 18296 7642 18352 7644
rect 18376 7642 18432 7644
rect 18456 7642 18512 7644
rect 18216 7590 18262 7642
rect 18262 7590 18272 7642
rect 18296 7590 18326 7642
rect 18326 7590 18338 7642
rect 18338 7590 18352 7642
rect 18376 7590 18390 7642
rect 18390 7590 18402 7642
rect 18402 7590 18432 7642
rect 18456 7590 18466 7642
rect 18466 7590 18512 7642
rect 18216 7588 18272 7590
rect 18296 7588 18352 7590
rect 18376 7588 18432 7590
rect 18456 7588 18512 7590
rect 1556 7098 1612 7100
rect 1636 7098 1692 7100
rect 1716 7098 1772 7100
rect 1796 7098 1852 7100
rect 1556 7046 1602 7098
rect 1602 7046 1612 7098
rect 1636 7046 1666 7098
rect 1666 7046 1678 7098
rect 1678 7046 1692 7098
rect 1716 7046 1730 7098
rect 1730 7046 1742 7098
rect 1742 7046 1772 7098
rect 1796 7046 1806 7098
rect 1806 7046 1852 7098
rect 1556 7044 1612 7046
rect 1636 7044 1692 7046
rect 1716 7044 1772 7046
rect 1796 7044 1852 7046
rect 5556 7098 5612 7100
rect 5636 7098 5692 7100
rect 5716 7098 5772 7100
rect 5796 7098 5852 7100
rect 5556 7046 5602 7098
rect 5602 7046 5612 7098
rect 5636 7046 5666 7098
rect 5666 7046 5678 7098
rect 5678 7046 5692 7098
rect 5716 7046 5730 7098
rect 5730 7046 5742 7098
rect 5742 7046 5772 7098
rect 5796 7046 5806 7098
rect 5806 7046 5852 7098
rect 5556 7044 5612 7046
rect 5636 7044 5692 7046
rect 5716 7044 5772 7046
rect 5796 7044 5852 7046
rect 9556 7098 9612 7100
rect 9636 7098 9692 7100
rect 9716 7098 9772 7100
rect 9796 7098 9852 7100
rect 9556 7046 9602 7098
rect 9602 7046 9612 7098
rect 9636 7046 9666 7098
rect 9666 7046 9678 7098
rect 9678 7046 9692 7098
rect 9716 7046 9730 7098
rect 9730 7046 9742 7098
rect 9742 7046 9772 7098
rect 9796 7046 9806 7098
rect 9806 7046 9852 7098
rect 9556 7044 9612 7046
rect 9636 7044 9692 7046
rect 9716 7044 9772 7046
rect 9796 7044 9852 7046
rect 13556 7098 13612 7100
rect 13636 7098 13692 7100
rect 13716 7098 13772 7100
rect 13796 7098 13852 7100
rect 13556 7046 13602 7098
rect 13602 7046 13612 7098
rect 13636 7046 13666 7098
rect 13666 7046 13678 7098
rect 13678 7046 13692 7098
rect 13716 7046 13730 7098
rect 13730 7046 13742 7098
rect 13742 7046 13772 7098
rect 13796 7046 13806 7098
rect 13806 7046 13852 7098
rect 13556 7044 13612 7046
rect 13636 7044 13692 7046
rect 13716 7044 13772 7046
rect 13796 7044 13852 7046
rect 17556 7098 17612 7100
rect 17636 7098 17692 7100
rect 17716 7098 17772 7100
rect 17796 7098 17852 7100
rect 17556 7046 17602 7098
rect 17602 7046 17612 7098
rect 17636 7046 17666 7098
rect 17666 7046 17678 7098
rect 17678 7046 17692 7098
rect 17716 7046 17730 7098
rect 17730 7046 17742 7098
rect 17742 7046 17772 7098
rect 17796 7046 17806 7098
rect 17806 7046 17852 7098
rect 17556 7044 17612 7046
rect 17636 7044 17692 7046
rect 17716 7044 17772 7046
rect 17796 7044 17852 7046
rect 2216 6554 2272 6556
rect 2296 6554 2352 6556
rect 2376 6554 2432 6556
rect 2456 6554 2512 6556
rect 2216 6502 2262 6554
rect 2262 6502 2272 6554
rect 2296 6502 2326 6554
rect 2326 6502 2338 6554
rect 2338 6502 2352 6554
rect 2376 6502 2390 6554
rect 2390 6502 2402 6554
rect 2402 6502 2432 6554
rect 2456 6502 2466 6554
rect 2466 6502 2512 6554
rect 2216 6500 2272 6502
rect 2296 6500 2352 6502
rect 2376 6500 2432 6502
rect 2456 6500 2512 6502
rect 6216 6554 6272 6556
rect 6296 6554 6352 6556
rect 6376 6554 6432 6556
rect 6456 6554 6512 6556
rect 6216 6502 6262 6554
rect 6262 6502 6272 6554
rect 6296 6502 6326 6554
rect 6326 6502 6338 6554
rect 6338 6502 6352 6554
rect 6376 6502 6390 6554
rect 6390 6502 6402 6554
rect 6402 6502 6432 6554
rect 6456 6502 6466 6554
rect 6466 6502 6512 6554
rect 6216 6500 6272 6502
rect 6296 6500 6352 6502
rect 6376 6500 6432 6502
rect 6456 6500 6512 6502
rect 10216 6554 10272 6556
rect 10296 6554 10352 6556
rect 10376 6554 10432 6556
rect 10456 6554 10512 6556
rect 10216 6502 10262 6554
rect 10262 6502 10272 6554
rect 10296 6502 10326 6554
rect 10326 6502 10338 6554
rect 10338 6502 10352 6554
rect 10376 6502 10390 6554
rect 10390 6502 10402 6554
rect 10402 6502 10432 6554
rect 10456 6502 10466 6554
rect 10466 6502 10512 6554
rect 10216 6500 10272 6502
rect 10296 6500 10352 6502
rect 10376 6500 10432 6502
rect 10456 6500 10512 6502
rect 14216 6554 14272 6556
rect 14296 6554 14352 6556
rect 14376 6554 14432 6556
rect 14456 6554 14512 6556
rect 14216 6502 14262 6554
rect 14262 6502 14272 6554
rect 14296 6502 14326 6554
rect 14326 6502 14338 6554
rect 14338 6502 14352 6554
rect 14376 6502 14390 6554
rect 14390 6502 14402 6554
rect 14402 6502 14432 6554
rect 14456 6502 14466 6554
rect 14466 6502 14512 6554
rect 14216 6500 14272 6502
rect 14296 6500 14352 6502
rect 14376 6500 14432 6502
rect 14456 6500 14512 6502
rect 18216 6554 18272 6556
rect 18296 6554 18352 6556
rect 18376 6554 18432 6556
rect 18456 6554 18512 6556
rect 18216 6502 18262 6554
rect 18262 6502 18272 6554
rect 18296 6502 18326 6554
rect 18326 6502 18338 6554
rect 18338 6502 18352 6554
rect 18376 6502 18390 6554
rect 18390 6502 18402 6554
rect 18402 6502 18432 6554
rect 18456 6502 18466 6554
rect 18466 6502 18512 6554
rect 18216 6500 18272 6502
rect 18296 6500 18352 6502
rect 18376 6500 18432 6502
rect 18456 6500 18512 6502
rect 1556 6010 1612 6012
rect 1636 6010 1692 6012
rect 1716 6010 1772 6012
rect 1796 6010 1852 6012
rect 1556 5958 1602 6010
rect 1602 5958 1612 6010
rect 1636 5958 1666 6010
rect 1666 5958 1678 6010
rect 1678 5958 1692 6010
rect 1716 5958 1730 6010
rect 1730 5958 1742 6010
rect 1742 5958 1772 6010
rect 1796 5958 1806 6010
rect 1806 5958 1852 6010
rect 1556 5956 1612 5958
rect 1636 5956 1692 5958
rect 1716 5956 1772 5958
rect 1796 5956 1852 5958
rect 5556 6010 5612 6012
rect 5636 6010 5692 6012
rect 5716 6010 5772 6012
rect 5796 6010 5852 6012
rect 5556 5958 5602 6010
rect 5602 5958 5612 6010
rect 5636 5958 5666 6010
rect 5666 5958 5678 6010
rect 5678 5958 5692 6010
rect 5716 5958 5730 6010
rect 5730 5958 5742 6010
rect 5742 5958 5772 6010
rect 5796 5958 5806 6010
rect 5806 5958 5852 6010
rect 5556 5956 5612 5958
rect 5636 5956 5692 5958
rect 5716 5956 5772 5958
rect 5796 5956 5852 5958
rect 9556 6010 9612 6012
rect 9636 6010 9692 6012
rect 9716 6010 9772 6012
rect 9796 6010 9852 6012
rect 9556 5958 9602 6010
rect 9602 5958 9612 6010
rect 9636 5958 9666 6010
rect 9666 5958 9678 6010
rect 9678 5958 9692 6010
rect 9716 5958 9730 6010
rect 9730 5958 9742 6010
rect 9742 5958 9772 6010
rect 9796 5958 9806 6010
rect 9806 5958 9852 6010
rect 9556 5956 9612 5958
rect 9636 5956 9692 5958
rect 9716 5956 9772 5958
rect 9796 5956 9852 5958
rect 13556 6010 13612 6012
rect 13636 6010 13692 6012
rect 13716 6010 13772 6012
rect 13796 6010 13852 6012
rect 13556 5958 13602 6010
rect 13602 5958 13612 6010
rect 13636 5958 13666 6010
rect 13666 5958 13678 6010
rect 13678 5958 13692 6010
rect 13716 5958 13730 6010
rect 13730 5958 13742 6010
rect 13742 5958 13772 6010
rect 13796 5958 13806 6010
rect 13806 5958 13852 6010
rect 13556 5956 13612 5958
rect 13636 5956 13692 5958
rect 13716 5956 13772 5958
rect 13796 5956 13852 5958
rect 17556 6010 17612 6012
rect 17636 6010 17692 6012
rect 17716 6010 17772 6012
rect 17796 6010 17852 6012
rect 17556 5958 17602 6010
rect 17602 5958 17612 6010
rect 17636 5958 17666 6010
rect 17666 5958 17678 6010
rect 17678 5958 17692 6010
rect 17716 5958 17730 6010
rect 17730 5958 17742 6010
rect 17742 5958 17772 6010
rect 17796 5958 17806 6010
rect 17806 5958 17852 6010
rect 17556 5956 17612 5958
rect 17636 5956 17692 5958
rect 17716 5956 17772 5958
rect 17796 5956 17852 5958
rect 2216 5466 2272 5468
rect 2296 5466 2352 5468
rect 2376 5466 2432 5468
rect 2456 5466 2512 5468
rect 2216 5414 2262 5466
rect 2262 5414 2272 5466
rect 2296 5414 2326 5466
rect 2326 5414 2338 5466
rect 2338 5414 2352 5466
rect 2376 5414 2390 5466
rect 2390 5414 2402 5466
rect 2402 5414 2432 5466
rect 2456 5414 2466 5466
rect 2466 5414 2512 5466
rect 2216 5412 2272 5414
rect 2296 5412 2352 5414
rect 2376 5412 2432 5414
rect 2456 5412 2512 5414
rect 6216 5466 6272 5468
rect 6296 5466 6352 5468
rect 6376 5466 6432 5468
rect 6456 5466 6512 5468
rect 6216 5414 6262 5466
rect 6262 5414 6272 5466
rect 6296 5414 6326 5466
rect 6326 5414 6338 5466
rect 6338 5414 6352 5466
rect 6376 5414 6390 5466
rect 6390 5414 6402 5466
rect 6402 5414 6432 5466
rect 6456 5414 6466 5466
rect 6466 5414 6512 5466
rect 6216 5412 6272 5414
rect 6296 5412 6352 5414
rect 6376 5412 6432 5414
rect 6456 5412 6512 5414
rect 10216 5466 10272 5468
rect 10296 5466 10352 5468
rect 10376 5466 10432 5468
rect 10456 5466 10512 5468
rect 10216 5414 10262 5466
rect 10262 5414 10272 5466
rect 10296 5414 10326 5466
rect 10326 5414 10338 5466
rect 10338 5414 10352 5466
rect 10376 5414 10390 5466
rect 10390 5414 10402 5466
rect 10402 5414 10432 5466
rect 10456 5414 10466 5466
rect 10466 5414 10512 5466
rect 10216 5412 10272 5414
rect 10296 5412 10352 5414
rect 10376 5412 10432 5414
rect 10456 5412 10512 5414
rect 14216 5466 14272 5468
rect 14296 5466 14352 5468
rect 14376 5466 14432 5468
rect 14456 5466 14512 5468
rect 14216 5414 14262 5466
rect 14262 5414 14272 5466
rect 14296 5414 14326 5466
rect 14326 5414 14338 5466
rect 14338 5414 14352 5466
rect 14376 5414 14390 5466
rect 14390 5414 14402 5466
rect 14402 5414 14432 5466
rect 14456 5414 14466 5466
rect 14466 5414 14512 5466
rect 14216 5412 14272 5414
rect 14296 5412 14352 5414
rect 14376 5412 14432 5414
rect 14456 5412 14512 5414
rect 18216 5466 18272 5468
rect 18296 5466 18352 5468
rect 18376 5466 18432 5468
rect 18456 5466 18512 5468
rect 18216 5414 18262 5466
rect 18262 5414 18272 5466
rect 18296 5414 18326 5466
rect 18326 5414 18338 5466
rect 18338 5414 18352 5466
rect 18376 5414 18390 5466
rect 18390 5414 18402 5466
rect 18402 5414 18432 5466
rect 18456 5414 18466 5466
rect 18466 5414 18512 5466
rect 18216 5412 18272 5414
rect 18296 5412 18352 5414
rect 18376 5412 18432 5414
rect 18456 5412 18512 5414
rect 1556 4922 1612 4924
rect 1636 4922 1692 4924
rect 1716 4922 1772 4924
rect 1796 4922 1852 4924
rect 1556 4870 1602 4922
rect 1602 4870 1612 4922
rect 1636 4870 1666 4922
rect 1666 4870 1678 4922
rect 1678 4870 1692 4922
rect 1716 4870 1730 4922
rect 1730 4870 1742 4922
rect 1742 4870 1772 4922
rect 1796 4870 1806 4922
rect 1806 4870 1852 4922
rect 1556 4868 1612 4870
rect 1636 4868 1692 4870
rect 1716 4868 1772 4870
rect 1796 4868 1852 4870
rect 5556 4922 5612 4924
rect 5636 4922 5692 4924
rect 5716 4922 5772 4924
rect 5796 4922 5852 4924
rect 5556 4870 5602 4922
rect 5602 4870 5612 4922
rect 5636 4870 5666 4922
rect 5666 4870 5678 4922
rect 5678 4870 5692 4922
rect 5716 4870 5730 4922
rect 5730 4870 5742 4922
rect 5742 4870 5772 4922
rect 5796 4870 5806 4922
rect 5806 4870 5852 4922
rect 5556 4868 5612 4870
rect 5636 4868 5692 4870
rect 5716 4868 5772 4870
rect 5796 4868 5852 4870
rect 9556 4922 9612 4924
rect 9636 4922 9692 4924
rect 9716 4922 9772 4924
rect 9796 4922 9852 4924
rect 9556 4870 9602 4922
rect 9602 4870 9612 4922
rect 9636 4870 9666 4922
rect 9666 4870 9678 4922
rect 9678 4870 9692 4922
rect 9716 4870 9730 4922
rect 9730 4870 9742 4922
rect 9742 4870 9772 4922
rect 9796 4870 9806 4922
rect 9806 4870 9852 4922
rect 9556 4868 9612 4870
rect 9636 4868 9692 4870
rect 9716 4868 9772 4870
rect 9796 4868 9852 4870
rect 13556 4922 13612 4924
rect 13636 4922 13692 4924
rect 13716 4922 13772 4924
rect 13796 4922 13852 4924
rect 13556 4870 13602 4922
rect 13602 4870 13612 4922
rect 13636 4870 13666 4922
rect 13666 4870 13678 4922
rect 13678 4870 13692 4922
rect 13716 4870 13730 4922
rect 13730 4870 13742 4922
rect 13742 4870 13772 4922
rect 13796 4870 13806 4922
rect 13806 4870 13852 4922
rect 13556 4868 13612 4870
rect 13636 4868 13692 4870
rect 13716 4868 13772 4870
rect 13796 4868 13852 4870
rect 17556 4922 17612 4924
rect 17636 4922 17692 4924
rect 17716 4922 17772 4924
rect 17796 4922 17852 4924
rect 17556 4870 17602 4922
rect 17602 4870 17612 4922
rect 17636 4870 17666 4922
rect 17666 4870 17678 4922
rect 17678 4870 17692 4922
rect 17716 4870 17730 4922
rect 17730 4870 17742 4922
rect 17742 4870 17772 4922
rect 17796 4870 17806 4922
rect 17806 4870 17852 4922
rect 17556 4868 17612 4870
rect 17636 4868 17692 4870
rect 17716 4868 17772 4870
rect 17796 4868 17852 4870
rect 2216 4378 2272 4380
rect 2296 4378 2352 4380
rect 2376 4378 2432 4380
rect 2456 4378 2512 4380
rect 2216 4326 2262 4378
rect 2262 4326 2272 4378
rect 2296 4326 2326 4378
rect 2326 4326 2338 4378
rect 2338 4326 2352 4378
rect 2376 4326 2390 4378
rect 2390 4326 2402 4378
rect 2402 4326 2432 4378
rect 2456 4326 2466 4378
rect 2466 4326 2512 4378
rect 2216 4324 2272 4326
rect 2296 4324 2352 4326
rect 2376 4324 2432 4326
rect 2456 4324 2512 4326
rect 6216 4378 6272 4380
rect 6296 4378 6352 4380
rect 6376 4378 6432 4380
rect 6456 4378 6512 4380
rect 6216 4326 6262 4378
rect 6262 4326 6272 4378
rect 6296 4326 6326 4378
rect 6326 4326 6338 4378
rect 6338 4326 6352 4378
rect 6376 4326 6390 4378
rect 6390 4326 6402 4378
rect 6402 4326 6432 4378
rect 6456 4326 6466 4378
rect 6466 4326 6512 4378
rect 6216 4324 6272 4326
rect 6296 4324 6352 4326
rect 6376 4324 6432 4326
rect 6456 4324 6512 4326
rect 10216 4378 10272 4380
rect 10296 4378 10352 4380
rect 10376 4378 10432 4380
rect 10456 4378 10512 4380
rect 10216 4326 10262 4378
rect 10262 4326 10272 4378
rect 10296 4326 10326 4378
rect 10326 4326 10338 4378
rect 10338 4326 10352 4378
rect 10376 4326 10390 4378
rect 10390 4326 10402 4378
rect 10402 4326 10432 4378
rect 10456 4326 10466 4378
rect 10466 4326 10512 4378
rect 10216 4324 10272 4326
rect 10296 4324 10352 4326
rect 10376 4324 10432 4326
rect 10456 4324 10512 4326
rect 14216 4378 14272 4380
rect 14296 4378 14352 4380
rect 14376 4378 14432 4380
rect 14456 4378 14512 4380
rect 14216 4326 14262 4378
rect 14262 4326 14272 4378
rect 14296 4326 14326 4378
rect 14326 4326 14338 4378
rect 14338 4326 14352 4378
rect 14376 4326 14390 4378
rect 14390 4326 14402 4378
rect 14402 4326 14432 4378
rect 14456 4326 14466 4378
rect 14466 4326 14512 4378
rect 14216 4324 14272 4326
rect 14296 4324 14352 4326
rect 14376 4324 14432 4326
rect 14456 4324 14512 4326
rect 18216 4378 18272 4380
rect 18296 4378 18352 4380
rect 18376 4378 18432 4380
rect 18456 4378 18512 4380
rect 18216 4326 18262 4378
rect 18262 4326 18272 4378
rect 18296 4326 18326 4378
rect 18326 4326 18338 4378
rect 18338 4326 18352 4378
rect 18376 4326 18390 4378
rect 18390 4326 18402 4378
rect 18402 4326 18432 4378
rect 18456 4326 18466 4378
rect 18466 4326 18512 4378
rect 18216 4324 18272 4326
rect 18296 4324 18352 4326
rect 18376 4324 18432 4326
rect 18456 4324 18512 4326
rect 1556 3834 1612 3836
rect 1636 3834 1692 3836
rect 1716 3834 1772 3836
rect 1796 3834 1852 3836
rect 1556 3782 1602 3834
rect 1602 3782 1612 3834
rect 1636 3782 1666 3834
rect 1666 3782 1678 3834
rect 1678 3782 1692 3834
rect 1716 3782 1730 3834
rect 1730 3782 1742 3834
rect 1742 3782 1772 3834
rect 1796 3782 1806 3834
rect 1806 3782 1852 3834
rect 1556 3780 1612 3782
rect 1636 3780 1692 3782
rect 1716 3780 1772 3782
rect 1796 3780 1852 3782
rect 5556 3834 5612 3836
rect 5636 3834 5692 3836
rect 5716 3834 5772 3836
rect 5796 3834 5852 3836
rect 5556 3782 5602 3834
rect 5602 3782 5612 3834
rect 5636 3782 5666 3834
rect 5666 3782 5678 3834
rect 5678 3782 5692 3834
rect 5716 3782 5730 3834
rect 5730 3782 5742 3834
rect 5742 3782 5772 3834
rect 5796 3782 5806 3834
rect 5806 3782 5852 3834
rect 5556 3780 5612 3782
rect 5636 3780 5692 3782
rect 5716 3780 5772 3782
rect 5796 3780 5852 3782
rect 9556 3834 9612 3836
rect 9636 3834 9692 3836
rect 9716 3834 9772 3836
rect 9796 3834 9852 3836
rect 9556 3782 9602 3834
rect 9602 3782 9612 3834
rect 9636 3782 9666 3834
rect 9666 3782 9678 3834
rect 9678 3782 9692 3834
rect 9716 3782 9730 3834
rect 9730 3782 9742 3834
rect 9742 3782 9772 3834
rect 9796 3782 9806 3834
rect 9806 3782 9852 3834
rect 9556 3780 9612 3782
rect 9636 3780 9692 3782
rect 9716 3780 9772 3782
rect 9796 3780 9852 3782
rect 13556 3834 13612 3836
rect 13636 3834 13692 3836
rect 13716 3834 13772 3836
rect 13796 3834 13852 3836
rect 13556 3782 13602 3834
rect 13602 3782 13612 3834
rect 13636 3782 13666 3834
rect 13666 3782 13678 3834
rect 13678 3782 13692 3834
rect 13716 3782 13730 3834
rect 13730 3782 13742 3834
rect 13742 3782 13772 3834
rect 13796 3782 13806 3834
rect 13806 3782 13852 3834
rect 13556 3780 13612 3782
rect 13636 3780 13692 3782
rect 13716 3780 13772 3782
rect 13796 3780 13852 3782
rect 17556 3834 17612 3836
rect 17636 3834 17692 3836
rect 17716 3834 17772 3836
rect 17796 3834 17852 3836
rect 17556 3782 17602 3834
rect 17602 3782 17612 3834
rect 17636 3782 17666 3834
rect 17666 3782 17678 3834
rect 17678 3782 17692 3834
rect 17716 3782 17730 3834
rect 17730 3782 17742 3834
rect 17742 3782 17772 3834
rect 17796 3782 17806 3834
rect 17806 3782 17852 3834
rect 17556 3780 17612 3782
rect 17636 3780 17692 3782
rect 17716 3780 17772 3782
rect 17796 3780 17852 3782
rect 2216 3290 2272 3292
rect 2296 3290 2352 3292
rect 2376 3290 2432 3292
rect 2456 3290 2512 3292
rect 2216 3238 2262 3290
rect 2262 3238 2272 3290
rect 2296 3238 2326 3290
rect 2326 3238 2338 3290
rect 2338 3238 2352 3290
rect 2376 3238 2390 3290
rect 2390 3238 2402 3290
rect 2402 3238 2432 3290
rect 2456 3238 2466 3290
rect 2466 3238 2512 3290
rect 2216 3236 2272 3238
rect 2296 3236 2352 3238
rect 2376 3236 2432 3238
rect 2456 3236 2512 3238
rect 6216 3290 6272 3292
rect 6296 3290 6352 3292
rect 6376 3290 6432 3292
rect 6456 3290 6512 3292
rect 6216 3238 6262 3290
rect 6262 3238 6272 3290
rect 6296 3238 6326 3290
rect 6326 3238 6338 3290
rect 6338 3238 6352 3290
rect 6376 3238 6390 3290
rect 6390 3238 6402 3290
rect 6402 3238 6432 3290
rect 6456 3238 6466 3290
rect 6466 3238 6512 3290
rect 6216 3236 6272 3238
rect 6296 3236 6352 3238
rect 6376 3236 6432 3238
rect 6456 3236 6512 3238
rect 10216 3290 10272 3292
rect 10296 3290 10352 3292
rect 10376 3290 10432 3292
rect 10456 3290 10512 3292
rect 10216 3238 10262 3290
rect 10262 3238 10272 3290
rect 10296 3238 10326 3290
rect 10326 3238 10338 3290
rect 10338 3238 10352 3290
rect 10376 3238 10390 3290
rect 10390 3238 10402 3290
rect 10402 3238 10432 3290
rect 10456 3238 10466 3290
rect 10466 3238 10512 3290
rect 10216 3236 10272 3238
rect 10296 3236 10352 3238
rect 10376 3236 10432 3238
rect 10456 3236 10512 3238
rect 14216 3290 14272 3292
rect 14296 3290 14352 3292
rect 14376 3290 14432 3292
rect 14456 3290 14512 3292
rect 14216 3238 14262 3290
rect 14262 3238 14272 3290
rect 14296 3238 14326 3290
rect 14326 3238 14338 3290
rect 14338 3238 14352 3290
rect 14376 3238 14390 3290
rect 14390 3238 14402 3290
rect 14402 3238 14432 3290
rect 14456 3238 14466 3290
rect 14466 3238 14512 3290
rect 14216 3236 14272 3238
rect 14296 3236 14352 3238
rect 14376 3236 14432 3238
rect 14456 3236 14512 3238
rect 18216 3290 18272 3292
rect 18296 3290 18352 3292
rect 18376 3290 18432 3292
rect 18456 3290 18512 3292
rect 18216 3238 18262 3290
rect 18262 3238 18272 3290
rect 18296 3238 18326 3290
rect 18326 3238 18338 3290
rect 18338 3238 18352 3290
rect 18376 3238 18390 3290
rect 18390 3238 18402 3290
rect 18402 3238 18432 3290
rect 18456 3238 18466 3290
rect 18466 3238 18512 3290
rect 18216 3236 18272 3238
rect 18296 3236 18352 3238
rect 18376 3236 18432 3238
rect 18456 3236 18512 3238
rect 1556 2746 1612 2748
rect 1636 2746 1692 2748
rect 1716 2746 1772 2748
rect 1796 2746 1852 2748
rect 1556 2694 1602 2746
rect 1602 2694 1612 2746
rect 1636 2694 1666 2746
rect 1666 2694 1678 2746
rect 1678 2694 1692 2746
rect 1716 2694 1730 2746
rect 1730 2694 1742 2746
rect 1742 2694 1772 2746
rect 1796 2694 1806 2746
rect 1806 2694 1852 2746
rect 1556 2692 1612 2694
rect 1636 2692 1692 2694
rect 1716 2692 1772 2694
rect 1796 2692 1852 2694
rect 5556 2746 5612 2748
rect 5636 2746 5692 2748
rect 5716 2746 5772 2748
rect 5796 2746 5852 2748
rect 5556 2694 5602 2746
rect 5602 2694 5612 2746
rect 5636 2694 5666 2746
rect 5666 2694 5678 2746
rect 5678 2694 5692 2746
rect 5716 2694 5730 2746
rect 5730 2694 5742 2746
rect 5742 2694 5772 2746
rect 5796 2694 5806 2746
rect 5806 2694 5852 2746
rect 5556 2692 5612 2694
rect 5636 2692 5692 2694
rect 5716 2692 5772 2694
rect 5796 2692 5852 2694
rect 9556 2746 9612 2748
rect 9636 2746 9692 2748
rect 9716 2746 9772 2748
rect 9796 2746 9852 2748
rect 9556 2694 9602 2746
rect 9602 2694 9612 2746
rect 9636 2694 9666 2746
rect 9666 2694 9678 2746
rect 9678 2694 9692 2746
rect 9716 2694 9730 2746
rect 9730 2694 9742 2746
rect 9742 2694 9772 2746
rect 9796 2694 9806 2746
rect 9806 2694 9852 2746
rect 9556 2692 9612 2694
rect 9636 2692 9692 2694
rect 9716 2692 9772 2694
rect 9796 2692 9852 2694
rect 13556 2746 13612 2748
rect 13636 2746 13692 2748
rect 13716 2746 13772 2748
rect 13796 2746 13852 2748
rect 13556 2694 13602 2746
rect 13602 2694 13612 2746
rect 13636 2694 13666 2746
rect 13666 2694 13678 2746
rect 13678 2694 13692 2746
rect 13716 2694 13730 2746
rect 13730 2694 13742 2746
rect 13742 2694 13772 2746
rect 13796 2694 13806 2746
rect 13806 2694 13852 2746
rect 13556 2692 13612 2694
rect 13636 2692 13692 2694
rect 13716 2692 13772 2694
rect 13796 2692 13852 2694
rect 17556 2746 17612 2748
rect 17636 2746 17692 2748
rect 17716 2746 17772 2748
rect 17796 2746 17852 2748
rect 17556 2694 17602 2746
rect 17602 2694 17612 2746
rect 17636 2694 17666 2746
rect 17666 2694 17678 2746
rect 17678 2694 17692 2746
rect 17716 2694 17730 2746
rect 17730 2694 17742 2746
rect 17742 2694 17772 2746
rect 17796 2694 17806 2746
rect 17806 2694 17852 2746
rect 17556 2692 17612 2694
rect 17636 2692 17692 2694
rect 17716 2692 17772 2694
rect 17796 2692 17852 2694
rect 2216 2202 2272 2204
rect 2296 2202 2352 2204
rect 2376 2202 2432 2204
rect 2456 2202 2512 2204
rect 2216 2150 2262 2202
rect 2262 2150 2272 2202
rect 2296 2150 2326 2202
rect 2326 2150 2338 2202
rect 2338 2150 2352 2202
rect 2376 2150 2390 2202
rect 2390 2150 2402 2202
rect 2402 2150 2432 2202
rect 2456 2150 2466 2202
rect 2466 2150 2512 2202
rect 2216 2148 2272 2150
rect 2296 2148 2352 2150
rect 2376 2148 2432 2150
rect 2456 2148 2512 2150
rect 6216 2202 6272 2204
rect 6296 2202 6352 2204
rect 6376 2202 6432 2204
rect 6456 2202 6512 2204
rect 6216 2150 6262 2202
rect 6262 2150 6272 2202
rect 6296 2150 6326 2202
rect 6326 2150 6338 2202
rect 6338 2150 6352 2202
rect 6376 2150 6390 2202
rect 6390 2150 6402 2202
rect 6402 2150 6432 2202
rect 6456 2150 6466 2202
rect 6466 2150 6512 2202
rect 6216 2148 6272 2150
rect 6296 2148 6352 2150
rect 6376 2148 6432 2150
rect 6456 2148 6512 2150
rect 10216 2202 10272 2204
rect 10296 2202 10352 2204
rect 10376 2202 10432 2204
rect 10456 2202 10512 2204
rect 10216 2150 10262 2202
rect 10262 2150 10272 2202
rect 10296 2150 10326 2202
rect 10326 2150 10338 2202
rect 10338 2150 10352 2202
rect 10376 2150 10390 2202
rect 10390 2150 10402 2202
rect 10402 2150 10432 2202
rect 10456 2150 10466 2202
rect 10466 2150 10512 2202
rect 10216 2148 10272 2150
rect 10296 2148 10352 2150
rect 10376 2148 10432 2150
rect 10456 2148 10512 2150
rect 14216 2202 14272 2204
rect 14296 2202 14352 2204
rect 14376 2202 14432 2204
rect 14456 2202 14512 2204
rect 14216 2150 14262 2202
rect 14262 2150 14272 2202
rect 14296 2150 14326 2202
rect 14326 2150 14338 2202
rect 14338 2150 14352 2202
rect 14376 2150 14390 2202
rect 14390 2150 14402 2202
rect 14402 2150 14432 2202
rect 14456 2150 14466 2202
rect 14466 2150 14512 2202
rect 14216 2148 14272 2150
rect 14296 2148 14352 2150
rect 14376 2148 14432 2150
rect 14456 2148 14512 2150
rect 18216 2202 18272 2204
rect 18296 2202 18352 2204
rect 18376 2202 18432 2204
rect 18456 2202 18512 2204
rect 18216 2150 18262 2202
rect 18262 2150 18272 2202
rect 18296 2150 18326 2202
rect 18326 2150 18338 2202
rect 18338 2150 18352 2202
rect 18376 2150 18390 2202
rect 18390 2150 18402 2202
rect 18402 2150 18432 2202
rect 18456 2150 18466 2202
rect 18466 2150 18512 2202
rect 18216 2148 18272 2150
rect 18296 2148 18352 2150
rect 18376 2148 18432 2150
rect 18456 2148 18512 2150
<< metal3 >>
rect 2206 17440 2522 17441
rect 2206 17376 2212 17440
rect 2276 17376 2292 17440
rect 2356 17376 2372 17440
rect 2436 17376 2452 17440
rect 2516 17376 2522 17440
rect 2206 17375 2522 17376
rect 6206 17440 6522 17441
rect 6206 17376 6212 17440
rect 6276 17376 6292 17440
rect 6356 17376 6372 17440
rect 6436 17376 6452 17440
rect 6516 17376 6522 17440
rect 6206 17375 6522 17376
rect 10206 17440 10522 17441
rect 10206 17376 10212 17440
rect 10276 17376 10292 17440
rect 10356 17376 10372 17440
rect 10436 17376 10452 17440
rect 10516 17376 10522 17440
rect 10206 17375 10522 17376
rect 14206 17440 14522 17441
rect 14206 17376 14212 17440
rect 14276 17376 14292 17440
rect 14356 17376 14372 17440
rect 14436 17376 14452 17440
rect 14516 17376 14522 17440
rect 14206 17375 14522 17376
rect 18206 17440 18522 17441
rect 18206 17376 18212 17440
rect 18276 17376 18292 17440
rect 18356 17376 18372 17440
rect 18436 17376 18452 17440
rect 18516 17376 18522 17440
rect 18206 17375 18522 17376
rect 1546 16896 1862 16897
rect 1546 16832 1552 16896
rect 1616 16832 1632 16896
rect 1696 16832 1712 16896
rect 1776 16832 1792 16896
rect 1856 16832 1862 16896
rect 1546 16831 1862 16832
rect 5546 16896 5862 16897
rect 5546 16832 5552 16896
rect 5616 16832 5632 16896
rect 5696 16832 5712 16896
rect 5776 16832 5792 16896
rect 5856 16832 5862 16896
rect 5546 16831 5862 16832
rect 9546 16896 9862 16897
rect 9546 16832 9552 16896
rect 9616 16832 9632 16896
rect 9696 16832 9712 16896
rect 9776 16832 9792 16896
rect 9856 16832 9862 16896
rect 9546 16831 9862 16832
rect 13546 16896 13862 16897
rect 13546 16832 13552 16896
rect 13616 16832 13632 16896
rect 13696 16832 13712 16896
rect 13776 16832 13792 16896
rect 13856 16832 13862 16896
rect 13546 16831 13862 16832
rect 17546 16896 17862 16897
rect 17546 16832 17552 16896
rect 17616 16832 17632 16896
rect 17696 16832 17712 16896
rect 17776 16832 17792 16896
rect 17856 16832 17862 16896
rect 17546 16831 17862 16832
rect 2206 16352 2522 16353
rect 2206 16288 2212 16352
rect 2276 16288 2292 16352
rect 2356 16288 2372 16352
rect 2436 16288 2452 16352
rect 2516 16288 2522 16352
rect 2206 16287 2522 16288
rect 6206 16352 6522 16353
rect 6206 16288 6212 16352
rect 6276 16288 6292 16352
rect 6356 16288 6372 16352
rect 6436 16288 6452 16352
rect 6516 16288 6522 16352
rect 6206 16287 6522 16288
rect 10206 16352 10522 16353
rect 10206 16288 10212 16352
rect 10276 16288 10292 16352
rect 10356 16288 10372 16352
rect 10436 16288 10452 16352
rect 10516 16288 10522 16352
rect 10206 16287 10522 16288
rect 14206 16352 14522 16353
rect 14206 16288 14212 16352
rect 14276 16288 14292 16352
rect 14356 16288 14372 16352
rect 14436 16288 14452 16352
rect 14516 16288 14522 16352
rect 14206 16287 14522 16288
rect 18206 16352 18522 16353
rect 18206 16288 18212 16352
rect 18276 16288 18292 16352
rect 18356 16288 18372 16352
rect 18436 16288 18452 16352
rect 18516 16288 18522 16352
rect 18206 16287 18522 16288
rect 1546 15808 1862 15809
rect 1546 15744 1552 15808
rect 1616 15744 1632 15808
rect 1696 15744 1712 15808
rect 1776 15744 1792 15808
rect 1856 15744 1862 15808
rect 1546 15743 1862 15744
rect 5546 15808 5862 15809
rect 5546 15744 5552 15808
rect 5616 15744 5632 15808
rect 5696 15744 5712 15808
rect 5776 15744 5792 15808
rect 5856 15744 5862 15808
rect 5546 15743 5862 15744
rect 9546 15808 9862 15809
rect 9546 15744 9552 15808
rect 9616 15744 9632 15808
rect 9696 15744 9712 15808
rect 9776 15744 9792 15808
rect 9856 15744 9862 15808
rect 9546 15743 9862 15744
rect 13546 15808 13862 15809
rect 13546 15744 13552 15808
rect 13616 15744 13632 15808
rect 13696 15744 13712 15808
rect 13776 15744 13792 15808
rect 13856 15744 13862 15808
rect 13546 15743 13862 15744
rect 17546 15808 17862 15809
rect 17546 15744 17552 15808
rect 17616 15744 17632 15808
rect 17696 15744 17712 15808
rect 17776 15744 17792 15808
rect 17856 15744 17862 15808
rect 17546 15743 17862 15744
rect 2206 15264 2522 15265
rect 2206 15200 2212 15264
rect 2276 15200 2292 15264
rect 2356 15200 2372 15264
rect 2436 15200 2452 15264
rect 2516 15200 2522 15264
rect 2206 15199 2522 15200
rect 6206 15264 6522 15265
rect 6206 15200 6212 15264
rect 6276 15200 6292 15264
rect 6356 15200 6372 15264
rect 6436 15200 6452 15264
rect 6516 15200 6522 15264
rect 6206 15199 6522 15200
rect 10206 15264 10522 15265
rect 10206 15200 10212 15264
rect 10276 15200 10292 15264
rect 10356 15200 10372 15264
rect 10436 15200 10452 15264
rect 10516 15200 10522 15264
rect 10206 15199 10522 15200
rect 14206 15264 14522 15265
rect 14206 15200 14212 15264
rect 14276 15200 14292 15264
rect 14356 15200 14372 15264
rect 14436 15200 14452 15264
rect 14516 15200 14522 15264
rect 14206 15199 14522 15200
rect 18206 15264 18522 15265
rect 18206 15200 18212 15264
rect 18276 15200 18292 15264
rect 18356 15200 18372 15264
rect 18436 15200 18452 15264
rect 18516 15200 18522 15264
rect 18206 15199 18522 15200
rect 1546 14720 1862 14721
rect 1546 14656 1552 14720
rect 1616 14656 1632 14720
rect 1696 14656 1712 14720
rect 1776 14656 1792 14720
rect 1856 14656 1862 14720
rect 1546 14655 1862 14656
rect 5546 14720 5862 14721
rect 5546 14656 5552 14720
rect 5616 14656 5632 14720
rect 5696 14656 5712 14720
rect 5776 14656 5792 14720
rect 5856 14656 5862 14720
rect 5546 14655 5862 14656
rect 9546 14720 9862 14721
rect 9546 14656 9552 14720
rect 9616 14656 9632 14720
rect 9696 14656 9712 14720
rect 9776 14656 9792 14720
rect 9856 14656 9862 14720
rect 9546 14655 9862 14656
rect 13546 14720 13862 14721
rect 13546 14656 13552 14720
rect 13616 14656 13632 14720
rect 13696 14656 13712 14720
rect 13776 14656 13792 14720
rect 13856 14656 13862 14720
rect 13546 14655 13862 14656
rect 17546 14720 17862 14721
rect 17546 14656 17552 14720
rect 17616 14656 17632 14720
rect 17696 14656 17712 14720
rect 17776 14656 17792 14720
rect 17856 14656 17862 14720
rect 17546 14655 17862 14656
rect 2206 14176 2522 14177
rect 2206 14112 2212 14176
rect 2276 14112 2292 14176
rect 2356 14112 2372 14176
rect 2436 14112 2452 14176
rect 2516 14112 2522 14176
rect 2206 14111 2522 14112
rect 6206 14176 6522 14177
rect 6206 14112 6212 14176
rect 6276 14112 6292 14176
rect 6356 14112 6372 14176
rect 6436 14112 6452 14176
rect 6516 14112 6522 14176
rect 6206 14111 6522 14112
rect 10206 14176 10522 14177
rect 10206 14112 10212 14176
rect 10276 14112 10292 14176
rect 10356 14112 10372 14176
rect 10436 14112 10452 14176
rect 10516 14112 10522 14176
rect 10206 14111 10522 14112
rect 14206 14176 14522 14177
rect 14206 14112 14212 14176
rect 14276 14112 14292 14176
rect 14356 14112 14372 14176
rect 14436 14112 14452 14176
rect 14516 14112 14522 14176
rect 14206 14111 14522 14112
rect 18206 14176 18522 14177
rect 18206 14112 18212 14176
rect 18276 14112 18292 14176
rect 18356 14112 18372 14176
rect 18436 14112 18452 14176
rect 18516 14112 18522 14176
rect 18206 14111 18522 14112
rect 1546 13632 1862 13633
rect 1546 13568 1552 13632
rect 1616 13568 1632 13632
rect 1696 13568 1712 13632
rect 1776 13568 1792 13632
rect 1856 13568 1862 13632
rect 1546 13567 1862 13568
rect 5546 13632 5862 13633
rect 5546 13568 5552 13632
rect 5616 13568 5632 13632
rect 5696 13568 5712 13632
rect 5776 13568 5792 13632
rect 5856 13568 5862 13632
rect 5546 13567 5862 13568
rect 9546 13632 9862 13633
rect 9546 13568 9552 13632
rect 9616 13568 9632 13632
rect 9696 13568 9712 13632
rect 9776 13568 9792 13632
rect 9856 13568 9862 13632
rect 9546 13567 9862 13568
rect 13546 13632 13862 13633
rect 13546 13568 13552 13632
rect 13616 13568 13632 13632
rect 13696 13568 13712 13632
rect 13776 13568 13792 13632
rect 13856 13568 13862 13632
rect 13546 13567 13862 13568
rect 17546 13632 17862 13633
rect 17546 13568 17552 13632
rect 17616 13568 17632 13632
rect 17696 13568 17712 13632
rect 17776 13568 17792 13632
rect 17856 13568 17862 13632
rect 17546 13567 17862 13568
rect 2206 13088 2522 13089
rect 2206 13024 2212 13088
rect 2276 13024 2292 13088
rect 2356 13024 2372 13088
rect 2436 13024 2452 13088
rect 2516 13024 2522 13088
rect 2206 13023 2522 13024
rect 6206 13088 6522 13089
rect 6206 13024 6212 13088
rect 6276 13024 6292 13088
rect 6356 13024 6372 13088
rect 6436 13024 6452 13088
rect 6516 13024 6522 13088
rect 6206 13023 6522 13024
rect 10206 13088 10522 13089
rect 10206 13024 10212 13088
rect 10276 13024 10292 13088
rect 10356 13024 10372 13088
rect 10436 13024 10452 13088
rect 10516 13024 10522 13088
rect 10206 13023 10522 13024
rect 14206 13088 14522 13089
rect 14206 13024 14212 13088
rect 14276 13024 14292 13088
rect 14356 13024 14372 13088
rect 14436 13024 14452 13088
rect 14516 13024 14522 13088
rect 14206 13023 14522 13024
rect 18206 13088 18522 13089
rect 18206 13024 18212 13088
rect 18276 13024 18292 13088
rect 18356 13024 18372 13088
rect 18436 13024 18452 13088
rect 18516 13024 18522 13088
rect 18206 13023 18522 13024
rect 1546 12544 1862 12545
rect 1546 12480 1552 12544
rect 1616 12480 1632 12544
rect 1696 12480 1712 12544
rect 1776 12480 1792 12544
rect 1856 12480 1862 12544
rect 1546 12479 1862 12480
rect 5546 12544 5862 12545
rect 5546 12480 5552 12544
rect 5616 12480 5632 12544
rect 5696 12480 5712 12544
rect 5776 12480 5792 12544
rect 5856 12480 5862 12544
rect 5546 12479 5862 12480
rect 9546 12544 9862 12545
rect 9546 12480 9552 12544
rect 9616 12480 9632 12544
rect 9696 12480 9712 12544
rect 9776 12480 9792 12544
rect 9856 12480 9862 12544
rect 9546 12479 9862 12480
rect 13546 12544 13862 12545
rect 13546 12480 13552 12544
rect 13616 12480 13632 12544
rect 13696 12480 13712 12544
rect 13776 12480 13792 12544
rect 13856 12480 13862 12544
rect 13546 12479 13862 12480
rect 17546 12544 17862 12545
rect 17546 12480 17552 12544
rect 17616 12480 17632 12544
rect 17696 12480 17712 12544
rect 17776 12480 17792 12544
rect 17856 12480 17862 12544
rect 17546 12479 17862 12480
rect 2206 12000 2522 12001
rect 2206 11936 2212 12000
rect 2276 11936 2292 12000
rect 2356 11936 2372 12000
rect 2436 11936 2452 12000
rect 2516 11936 2522 12000
rect 2206 11935 2522 11936
rect 6206 12000 6522 12001
rect 6206 11936 6212 12000
rect 6276 11936 6292 12000
rect 6356 11936 6372 12000
rect 6436 11936 6452 12000
rect 6516 11936 6522 12000
rect 6206 11935 6522 11936
rect 10206 12000 10522 12001
rect 10206 11936 10212 12000
rect 10276 11936 10292 12000
rect 10356 11936 10372 12000
rect 10436 11936 10452 12000
rect 10516 11936 10522 12000
rect 10206 11935 10522 11936
rect 14206 12000 14522 12001
rect 14206 11936 14212 12000
rect 14276 11936 14292 12000
rect 14356 11936 14372 12000
rect 14436 11936 14452 12000
rect 14516 11936 14522 12000
rect 14206 11935 14522 11936
rect 18206 12000 18522 12001
rect 18206 11936 18212 12000
rect 18276 11936 18292 12000
rect 18356 11936 18372 12000
rect 18436 11936 18452 12000
rect 18516 11936 18522 12000
rect 18206 11935 18522 11936
rect 841 11794 907 11797
rect 798 11792 907 11794
rect 798 11736 846 11792
rect 902 11736 907 11792
rect 798 11731 907 11736
rect 798 11688 858 11731
rect 0 11598 858 11688
rect 0 11568 800 11598
rect 1546 11456 1862 11457
rect 1546 11392 1552 11456
rect 1616 11392 1632 11456
rect 1696 11392 1712 11456
rect 1776 11392 1792 11456
rect 1856 11392 1862 11456
rect 1546 11391 1862 11392
rect 5546 11456 5862 11457
rect 5546 11392 5552 11456
rect 5616 11392 5632 11456
rect 5696 11392 5712 11456
rect 5776 11392 5792 11456
rect 5856 11392 5862 11456
rect 5546 11391 5862 11392
rect 9546 11456 9862 11457
rect 9546 11392 9552 11456
rect 9616 11392 9632 11456
rect 9696 11392 9712 11456
rect 9776 11392 9792 11456
rect 9856 11392 9862 11456
rect 9546 11391 9862 11392
rect 13546 11456 13862 11457
rect 13546 11392 13552 11456
rect 13616 11392 13632 11456
rect 13696 11392 13712 11456
rect 13776 11392 13792 11456
rect 13856 11392 13862 11456
rect 13546 11391 13862 11392
rect 17546 11456 17862 11457
rect 17546 11392 17552 11456
rect 17616 11392 17632 11456
rect 17696 11392 17712 11456
rect 17776 11392 17792 11456
rect 17856 11392 17862 11456
rect 17546 11391 17862 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 2206 10912 2522 10913
rect 2206 10848 2212 10912
rect 2276 10848 2292 10912
rect 2356 10848 2372 10912
rect 2436 10848 2452 10912
rect 2516 10848 2522 10912
rect 2206 10847 2522 10848
rect 6206 10912 6522 10913
rect 6206 10848 6212 10912
rect 6276 10848 6292 10912
rect 6356 10848 6372 10912
rect 6436 10848 6452 10912
rect 6516 10848 6522 10912
rect 6206 10847 6522 10848
rect 10206 10912 10522 10913
rect 10206 10848 10212 10912
rect 10276 10848 10292 10912
rect 10356 10848 10372 10912
rect 10436 10848 10452 10912
rect 10516 10848 10522 10912
rect 10206 10847 10522 10848
rect 14206 10912 14522 10913
rect 14206 10848 14212 10912
rect 14276 10848 14292 10912
rect 14356 10848 14372 10912
rect 14436 10848 14452 10912
rect 14516 10848 14522 10912
rect 14206 10847 14522 10848
rect 18206 10912 18522 10913
rect 18206 10848 18212 10912
rect 18276 10848 18292 10912
rect 18356 10848 18372 10912
rect 18436 10848 18452 10912
rect 18516 10848 18522 10912
rect 18206 10847 18522 10848
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 1546 10368 1862 10369
rect 1546 10304 1552 10368
rect 1616 10304 1632 10368
rect 1696 10304 1712 10368
rect 1776 10304 1792 10368
rect 1856 10304 1862 10368
rect 1546 10303 1862 10304
rect 5546 10368 5862 10369
rect 5546 10304 5552 10368
rect 5616 10304 5632 10368
rect 5696 10304 5712 10368
rect 5776 10304 5792 10368
rect 5856 10304 5862 10368
rect 5546 10303 5862 10304
rect 9546 10368 9862 10369
rect 9546 10304 9552 10368
rect 9616 10304 9632 10368
rect 9696 10304 9712 10368
rect 9776 10304 9792 10368
rect 9856 10304 9862 10368
rect 9546 10303 9862 10304
rect 13546 10368 13862 10369
rect 13546 10304 13552 10368
rect 13616 10304 13632 10368
rect 13696 10304 13712 10368
rect 13776 10304 13792 10368
rect 13856 10304 13862 10368
rect 13546 10303 13862 10304
rect 17546 10368 17862 10369
rect 17546 10304 17552 10368
rect 17616 10304 17632 10368
rect 17696 10304 17712 10368
rect 17776 10304 17792 10368
rect 17856 10304 17862 10368
rect 17546 10303 17862 10304
rect 18505 10298 18571 10301
rect 19200 10298 20000 10328
rect 18505 10296 20000 10298
rect 18505 10240 18510 10296
rect 18566 10240 20000 10296
rect 18505 10238 20000 10240
rect 0 10208 800 10238
rect 18505 10235 18571 10238
rect 19200 10208 20000 10238
rect 2206 9824 2522 9825
rect 2206 9760 2212 9824
rect 2276 9760 2292 9824
rect 2356 9760 2372 9824
rect 2436 9760 2452 9824
rect 2516 9760 2522 9824
rect 2206 9759 2522 9760
rect 6206 9824 6522 9825
rect 6206 9760 6212 9824
rect 6276 9760 6292 9824
rect 6356 9760 6372 9824
rect 6436 9760 6452 9824
rect 6516 9760 6522 9824
rect 6206 9759 6522 9760
rect 10206 9824 10522 9825
rect 10206 9760 10212 9824
rect 10276 9760 10292 9824
rect 10356 9760 10372 9824
rect 10436 9760 10452 9824
rect 10516 9760 10522 9824
rect 10206 9759 10522 9760
rect 14206 9824 14522 9825
rect 14206 9760 14212 9824
rect 14276 9760 14292 9824
rect 14356 9760 14372 9824
rect 14436 9760 14452 9824
rect 14516 9760 14522 9824
rect 14206 9759 14522 9760
rect 18206 9824 18522 9825
rect 18206 9760 18212 9824
rect 18276 9760 18292 9824
rect 18356 9760 18372 9824
rect 18436 9760 18452 9824
rect 18516 9760 18522 9824
rect 18206 9759 18522 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 1546 9280 1862 9281
rect 1546 9216 1552 9280
rect 1616 9216 1632 9280
rect 1696 9216 1712 9280
rect 1776 9216 1792 9280
rect 1856 9216 1862 9280
rect 1546 9215 1862 9216
rect 5546 9280 5862 9281
rect 5546 9216 5552 9280
rect 5616 9216 5632 9280
rect 5696 9216 5712 9280
rect 5776 9216 5792 9280
rect 5856 9216 5862 9280
rect 5546 9215 5862 9216
rect 9546 9280 9862 9281
rect 9546 9216 9552 9280
rect 9616 9216 9632 9280
rect 9696 9216 9712 9280
rect 9776 9216 9792 9280
rect 9856 9216 9862 9280
rect 9546 9215 9862 9216
rect 13546 9280 13862 9281
rect 13546 9216 13552 9280
rect 13616 9216 13632 9280
rect 13696 9216 13712 9280
rect 13776 9216 13792 9280
rect 13856 9216 13862 9280
rect 13546 9215 13862 9216
rect 17546 9280 17862 9281
rect 17546 9216 17552 9280
rect 17616 9216 17632 9280
rect 17696 9216 17712 9280
rect 17776 9216 17792 9280
rect 17856 9216 17862 9280
rect 17546 9215 17862 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 0 8848 800 8878
rect 2206 8736 2522 8737
rect 2206 8672 2212 8736
rect 2276 8672 2292 8736
rect 2356 8672 2372 8736
rect 2436 8672 2452 8736
rect 2516 8672 2522 8736
rect 2206 8671 2522 8672
rect 6206 8736 6522 8737
rect 6206 8672 6212 8736
rect 6276 8672 6292 8736
rect 6356 8672 6372 8736
rect 6436 8672 6452 8736
rect 6516 8672 6522 8736
rect 6206 8671 6522 8672
rect 10206 8736 10522 8737
rect 10206 8672 10212 8736
rect 10276 8672 10292 8736
rect 10356 8672 10372 8736
rect 10436 8672 10452 8736
rect 10516 8672 10522 8736
rect 10206 8671 10522 8672
rect 14206 8736 14522 8737
rect 14206 8672 14212 8736
rect 14276 8672 14292 8736
rect 14356 8672 14372 8736
rect 14436 8672 14452 8736
rect 14516 8672 14522 8736
rect 14206 8671 14522 8672
rect 18206 8736 18522 8737
rect 18206 8672 18212 8736
rect 18276 8672 18292 8736
rect 18356 8672 18372 8736
rect 18436 8672 18452 8736
rect 18516 8672 18522 8736
rect 18206 8671 18522 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 1546 8192 1862 8193
rect 1546 8128 1552 8192
rect 1616 8128 1632 8192
rect 1696 8128 1712 8192
rect 1776 8128 1792 8192
rect 1856 8128 1862 8192
rect 1546 8127 1862 8128
rect 5546 8192 5862 8193
rect 5546 8128 5552 8192
rect 5616 8128 5632 8192
rect 5696 8128 5712 8192
rect 5776 8128 5792 8192
rect 5856 8128 5862 8192
rect 5546 8127 5862 8128
rect 9546 8192 9862 8193
rect 9546 8128 9552 8192
rect 9616 8128 9632 8192
rect 9696 8128 9712 8192
rect 9776 8128 9792 8192
rect 9856 8128 9862 8192
rect 9546 8127 9862 8128
rect 13546 8192 13862 8193
rect 13546 8128 13552 8192
rect 13616 8128 13632 8192
rect 13696 8128 13712 8192
rect 13776 8128 13792 8192
rect 13856 8128 13862 8192
rect 13546 8127 13862 8128
rect 17546 8192 17862 8193
rect 17546 8128 17552 8192
rect 17616 8128 17632 8192
rect 17696 8128 17712 8192
rect 17776 8128 17792 8192
rect 17856 8128 17862 8192
rect 17546 8127 17862 8128
rect 2206 7648 2522 7649
rect 2206 7584 2212 7648
rect 2276 7584 2292 7648
rect 2356 7584 2372 7648
rect 2436 7584 2452 7648
rect 2516 7584 2522 7648
rect 2206 7583 2522 7584
rect 6206 7648 6522 7649
rect 6206 7584 6212 7648
rect 6276 7584 6292 7648
rect 6356 7584 6372 7648
rect 6436 7584 6452 7648
rect 6516 7584 6522 7648
rect 6206 7583 6522 7584
rect 10206 7648 10522 7649
rect 10206 7584 10212 7648
rect 10276 7584 10292 7648
rect 10356 7584 10372 7648
rect 10436 7584 10452 7648
rect 10516 7584 10522 7648
rect 10206 7583 10522 7584
rect 14206 7648 14522 7649
rect 14206 7584 14212 7648
rect 14276 7584 14292 7648
rect 14356 7584 14372 7648
rect 14436 7584 14452 7648
rect 14516 7584 14522 7648
rect 14206 7583 14522 7584
rect 18206 7648 18522 7649
rect 18206 7584 18212 7648
rect 18276 7584 18292 7648
rect 18356 7584 18372 7648
rect 18436 7584 18452 7648
rect 18516 7584 18522 7648
rect 18206 7583 18522 7584
rect 1546 7104 1862 7105
rect 1546 7040 1552 7104
rect 1616 7040 1632 7104
rect 1696 7040 1712 7104
rect 1776 7040 1792 7104
rect 1856 7040 1862 7104
rect 1546 7039 1862 7040
rect 5546 7104 5862 7105
rect 5546 7040 5552 7104
rect 5616 7040 5632 7104
rect 5696 7040 5712 7104
rect 5776 7040 5792 7104
rect 5856 7040 5862 7104
rect 5546 7039 5862 7040
rect 9546 7104 9862 7105
rect 9546 7040 9552 7104
rect 9616 7040 9632 7104
rect 9696 7040 9712 7104
rect 9776 7040 9792 7104
rect 9856 7040 9862 7104
rect 9546 7039 9862 7040
rect 13546 7104 13862 7105
rect 13546 7040 13552 7104
rect 13616 7040 13632 7104
rect 13696 7040 13712 7104
rect 13776 7040 13792 7104
rect 13856 7040 13862 7104
rect 13546 7039 13862 7040
rect 17546 7104 17862 7105
rect 17546 7040 17552 7104
rect 17616 7040 17632 7104
rect 17696 7040 17712 7104
rect 17776 7040 17792 7104
rect 17856 7040 17862 7104
rect 17546 7039 17862 7040
rect 2206 6560 2522 6561
rect 2206 6496 2212 6560
rect 2276 6496 2292 6560
rect 2356 6496 2372 6560
rect 2436 6496 2452 6560
rect 2516 6496 2522 6560
rect 2206 6495 2522 6496
rect 6206 6560 6522 6561
rect 6206 6496 6212 6560
rect 6276 6496 6292 6560
rect 6356 6496 6372 6560
rect 6436 6496 6452 6560
rect 6516 6496 6522 6560
rect 6206 6495 6522 6496
rect 10206 6560 10522 6561
rect 10206 6496 10212 6560
rect 10276 6496 10292 6560
rect 10356 6496 10372 6560
rect 10436 6496 10452 6560
rect 10516 6496 10522 6560
rect 10206 6495 10522 6496
rect 14206 6560 14522 6561
rect 14206 6496 14212 6560
rect 14276 6496 14292 6560
rect 14356 6496 14372 6560
rect 14436 6496 14452 6560
rect 14516 6496 14522 6560
rect 14206 6495 14522 6496
rect 18206 6560 18522 6561
rect 18206 6496 18212 6560
rect 18276 6496 18292 6560
rect 18356 6496 18372 6560
rect 18436 6496 18452 6560
rect 18516 6496 18522 6560
rect 18206 6495 18522 6496
rect 1546 6016 1862 6017
rect 1546 5952 1552 6016
rect 1616 5952 1632 6016
rect 1696 5952 1712 6016
rect 1776 5952 1792 6016
rect 1856 5952 1862 6016
rect 1546 5951 1862 5952
rect 5546 6016 5862 6017
rect 5546 5952 5552 6016
rect 5616 5952 5632 6016
rect 5696 5952 5712 6016
rect 5776 5952 5792 6016
rect 5856 5952 5862 6016
rect 5546 5951 5862 5952
rect 9546 6016 9862 6017
rect 9546 5952 9552 6016
rect 9616 5952 9632 6016
rect 9696 5952 9712 6016
rect 9776 5952 9792 6016
rect 9856 5952 9862 6016
rect 9546 5951 9862 5952
rect 13546 6016 13862 6017
rect 13546 5952 13552 6016
rect 13616 5952 13632 6016
rect 13696 5952 13712 6016
rect 13776 5952 13792 6016
rect 13856 5952 13862 6016
rect 13546 5951 13862 5952
rect 17546 6016 17862 6017
rect 17546 5952 17552 6016
rect 17616 5952 17632 6016
rect 17696 5952 17712 6016
rect 17776 5952 17792 6016
rect 17856 5952 17862 6016
rect 17546 5951 17862 5952
rect 2206 5472 2522 5473
rect 2206 5408 2212 5472
rect 2276 5408 2292 5472
rect 2356 5408 2372 5472
rect 2436 5408 2452 5472
rect 2516 5408 2522 5472
rect 2206 5407 2522 5408
rect 6206 5472 6522 5473
rect 6206 5408 6212 5472
rect 6276 5408 6292 5472
rect 6356 5408 6372 5472
rect 6436 5408 6452 5472
rect 6516 5408 6522 5472
rect 6206 5407 6522 5408
rect 10206 5472 10522 5473
rect 10206 5408 10212 5472
rect 10276 5408 10292 5472
rect 10356 5408 10372 5472
rect 10436 5408 10452 5472
rect 10516 5408 10522 5472
rect 10206 5407 10522 5408
rect 14206 5472 14522 5473
rect 14206 5408 14212 5472
rect 14276 5408 14292 5472
rect 14356 5408 14372 5472
rect 14436 5408 14452 5472
rect 14516 5408 14522 5472
rect 14206 5407 14522 5408
rect 18206 5472 18522 5473
rect 18206 5408 18212 5472
rect 18276 5408 18292 5472
rect 18356 5408 18372 5472
rect 18436 5408 18452 5472
rect 18516 5408 18522 5472
rect 18206 5407 18522 5408
rect 1546 4928 1862 4929
rect 1546 4864 1552 4928
rect 1616 4864 1632 4928
rect 1696 4864 1712 4928
rect 1776 4864 1792 4928
rect 1856 4864 1862 4928
rect 1546 4863 1862 4864
rect 5546 4928 5862 4929
rect 5546 4864 5552 4928
rect 5616 4864 5632 4928
rect 5696 4864 5712 4928
rect 5776 4864 5792 4928
rect 5856 4864 5862 4928
rect 5546 4863 5862 4864
rect 9546 4928 9862 4929
rect 9546 4864 9552 4928
rect 9616 4864 9632 4928
rect 9696 4864 9712 4928
rect 9776 4864 9792 4928
rect 9856 4864 9862 4928
rect 9546 4863 9862 4864
rect 13546 4928 13862 4929
rect 13546 4864 13552 4928
rect 13616 4864 13632 4928
rect 13696 4864 13712 4928
rect 13776 4864 13792 4928
rect 13856 4864 13862 4928
rect 13546 4863 13862 4864
rect 17546 4928 17862 4929
rect 17546 4864 17552 4928
rect 17616 4864 17632 4928
rect 17696 4864 17712 4928
rect 17776 4864 17792 4928
rect 17856 4864 17862 4928
rect 17546 4863 17862 4864
rect 2206 4384 2522 4385
rect 2206 4320 2212 4384
rect 2276 4320 2292 4384
rect 2356 4320 2372 4384
rect 2436 4320 2452 4384
rect 2516 4320 2522 4384
rect 2206 4319 2522 4320
rect 6206 4384 6522 4385
rect 6206 4320 6212 4384
rect 6276 4320 6292 4384
rect 6356 4320 6372 4384
rect 6436 4320 6452 4384
rect 6516 4320 6522 4384
rect 6206 4319 6522 4320
rect 10206 4384 10522 4385
rect 10206 4320 10212 4384
rect 10276 4320 10292 4384
rect 10356 4320 10372 4384
rect 10436 4320 10452 4384
rect 10516 4320 10522 4384
rect 10206 4319 10522 4320
rect 14206 4384 14522 4385
rect 14206 4320 14212 4384
rect 14276 4320 14292 4384
rect 14356 4320 14372 4384
rect 14436 4320 14452 4384
rect 14516 4320 14522 4384
rect 14206 4319 14522 4320
rect 18206 4384 18522 4385
rect 18206 4320 18212 4384
rect 18276 4320 18292 4384
rect 18356 4320 18372 4384
rect 18436 4320 18452 4384
rect 18516 4320 18522 4384
rect 18206 4319 18522 4320
rect 1546 3840 1862 3841
rect 1546 3776 1552 3840
rect 1616 3776 1632 3840
rect 1696 3776 1712 3840
rect 1776 3776 1792 3840
rect 1856 3776 1862 3840
rect 1546 3775 1862 3776
rect 5546 3840 5862 3841
rect 5546 3776 5552 3840
rect 5616 3776 5632 3840
rect 5696 3776 5712 3840
rect 5776 3776 5792 3840
rect 5856 3776 5862 3840
rect 5546 3775 5862 3776
rect 9546 3840 9862 3841
rect 9546 3776 9552 3840
rect 9616 3776 9632 3840
rect 9696 3776 9712 3840
rect 9776 3776 9792 3840
rect 9856 3776 9862 3840
rect 9546 3775 9862 3776
rect 13546 3840 13862 3841
rect 13546 3776 13552 3840
rect 13616 3776 13632 3840
rect 13696 3776 13712 3840
rect 13776 3776 13792 3840
rect 13856 3776 13862 3840
rect 13546 3775 13862 3776
rect 17546 3840 17862 3841
rect 17546 3776 17552 3840
rect 17616 3776 17632 3840
rect 17696 3776 17712 3840
rect 17776 3776 17792 3840
rect 17856 3776 17862 3840
rect 17546 3775 17862 3776
rect 2206 3296 2522 3297
rect 2206 3232 2212 3296
rect 2276 3232 2292 3296
rect 2356 3232 2372 3296
rect 2436 3232 2452 3296
rect 2516 3232 2522 3296
rect 2206 3231 2522 3232
rect 6206 3296 6522 3297
rect 6206 3232 6212 3296
rect 6276 3232 6292 3296
rect 6356 3232 6372 3296
rect 6436 3232 6452 3296
rect 6516 3232 6522 3296
rect 6206 3231 6522 3232
rect 10206 3296 10522 3297
rect 10206 3232 10212 3296
rect 10276 3232 10292 3296
rect 10356 3232 10372 3296
rect 10436 3232 10452 3296
rect 10516 3232 10522 3296
rect 10206 3231 10522 3232
rect 14206 3296 14522 3297
rect 14206 3232 14212 3296
rect 14276 3232 14292 3296
rect 14356 3232 14372 3296
rect 14436 3232 14452 3296
rect 14516 3232 14522 3296
rect 14206 3231 14522 3232
rect 18206 3296 18522 3297
rect 18206 3232 18212 3296
rect 18276 3232 18292 3296
rect 18356 3232 18372 3296
rect 18436 3232 18452 3296
rect 18516 3232 18522 3296
rect 18206 3231 18522 3232
rect 1546 2752 1862 2753
rect 1546 2688 1552 2752
rect 1616 2688 1632 2752
rect 1696 2688 1712 2752
rect 1776 2688 1792 2752
rect 1856 2688 1862 2752
rect 1546 2687 1862 2688
rect 5546 2752 5862 2753
rect 5546 2688 5552 2752
rect 5616 2688 5632 2752
rect 5696 2688 5712 2752
rect 5776 2688 5792 2752
rect 5856 2688 5862 2752
rect 5546 2687 5862 2688
rect 9546 2752 9862 2753
rect 9546 2688 9552 2752
rect 9616 2688 9632 2752
rect 9696 2688 9712 2752
rect 9776 2688 9792 2752
rect 9856 2688 9862 2752
rect 9546 2687 9862 2688
rect 13546 2752 13862 2753
rect 13546 2688 13552 2752
rect 13616 2688 13632 2752
rect 13696 2688 13712 2752
rect 13776 2688 13792 2752
rect 13856 2688 13862 2752
rect 13546 2687 13862 2688
rect 17546 2752 17862 2753
rect 17546 2688 17552 2752
rect 17616 2688 17632 2752
rect 17696 2688 17712 2752
rect 17776 2688 17792 2752
rect 17856 2688 17862 2752
rect 17546 2687 17862 2688
rect 2206 2208 2522 2209
rect 2206 2144 2212 2208
rect 2276 2144 2292 2208
rect 2356 2144 2372 2208
rect 2436 2144 2452 2208
rect 2516 2144 2522 2208
rect 2206 2143 2522 2144
rect 6206 2208 6522 2209
rect 6206 2144 6212 2208
rect 6276 2144 6292 2208
rect 6356 2144 6372 2208
rect 6436 2144 6452 2208
rect 6516 2144 6522 2208
rect 6206 2143 6522 2144
rect 10206 2208 10522 2209
rect 10206 2144 10212 2208
rect 10276 2144 10292 2208
rect 10356 2144 10372 2208
rect 10436 2144 10452 2208
rect 10516 2144 10522 2208
rect 10206 2143 10522 2144
rect 14206 2208 14522 2209
rect 14206 2144 14212 2208
rect 14276 2144 14292 2208
rect 14356 2144 14372 2208
rect 14436 2144 14452 2208
rect 14516 2144 14522 2208
rect 14206 2143 14522 2144
rect 18206 2208 18522 2209
rect 18206 2144 18212 2208
rect 18276 2144 18292 2208
rect 18356 2144 18372 2208
rect 18436 2144 18452 2208
rect 18516 2144 18522 2208
rect 18206 2143 18522 2144
<< via3 >>
rect 2212 17436 2276 17440
rect 2212 17380 2216 17436
rect 2216 17380 2272 17436
rect 2272 17380 2276 17436
rect 2212 17376 2276 17380
rect 2292 17436 2356 17440
rect 2292 17380 2296 17436
rect 2296 17380 2352 17436
rect 2352 17380 2356 17436
rect 2292 17376 2356 17380
rect 2372 17436 2436 17440
rect 2372 17380 2376 17436
rect 2376 17380 2432 17436
rect 2432 17380 2436 17436
rect 2372 17376 2436 17380
rect 2452 17436 2516 17440
rect 2452 17380 2456 17436
rect 2456 17380 2512 17436
rect 2512 17380 2516 17436
rect 2452 17376 2516 17380
rect 6212 17436 6276 17440
rect 6212 17380 6216 17436
rect 6216 17380 6272 17436
rect 6272 17380 6276 17436
rect 6212 17376 6276 17380
rect 6292 17436 6356 17440
rect 6292 17380 6296 17436
rect 6296 17380 6352 17436
rect 6352 17380 6356 17436
rect 6292 17376 6356 17380
rect 6372 17436 6436 17440
rect 6372 17380 6376 17436
rect 6376 17380 6432 17436
rect 6432 17380 6436 17436
rect 6372 17376 6436 17380
rect 6452 17436 6516 17440
rect 6452 17380 6456 17436
rect 6456 17380 6512 17436
rect 6512 17380 6516 17436
rect 6452 17376 6516 17380
rect 10212 17436 10276 17440
rect 10212 17380 10216 17436
rect 10216 17380 10272 17436
rect 10272 17380 10276 17436
rect 10212 17376 10276 17380
rect 10292 17436 10356 17440
rect 10292 17380 10296 17436
rect 10296 17380 10352 17436
rect 10352 17380 10356 17436
rect 10292 17376 10356 17380
rect 10372 17436 10436 17440
rect 10372 17380 10376 17436
rect 10376 17380 10432 17436
rect 10432 17380 10436 17436
rect 10372 17376 10436 17380
rect 10452 17436 10516 17440
rect 10452 17380 10456 17436
rect 10456 17380 10512 17436
rect 10512 17380 10516 17436
rect 10452 17376 10516 17380
rect 14212 17436 14276 17440
rect 14212 17380 14216 17436
rect 14216 17380 14272 17436
rect 14272 17380 14276 17436
rect 14212 17376 14276 17380
rect 14292 17436 14356 17440
rect 14292 17380 14296 17436
rect 14296 17380 14352 17436
rect 14352 17380 14356 17436
rect 14292 17376 14356 17380
rect 14372 17436 14436 17440
rect 14372 17380 14376 17436
rect 14376 17380 14432 17436
rect 14432 17380 14436 17436
rect 14372 17376 14436 17380
rect 14452 17436 14516 17440
rect 14452 17380 14456 17436
rect 14456 17380 14512 17436
rect 14512 17380 14516 17436
rect 14452 17376 14516 17380
rect 18212 17436 18276 17440
rect 18212 17380 18216 17436
rect 18216 17380 18272 17436
rect 18272 17380 18276 17436
rect 18212 17376 18276 17380
rect 18292 17436 18356 17440
rect 18292 17380 18296 17436
rect 18296 17380 18352 17436
rect 18352 17380 18356 17436
rect 18292 17376 18356 17380
rect 18372 17436 18436 17440
rect 18372 17380 18376 17436
rect 18376 17380 18432 17436
rect 18432 17380 18436 17436
rect 18372 17376 18436 17380
rect 18452 17436 18516 17440
rect 18452 17380 18456 17436
rect 18456 17380 18512 17436
rect 18512 17380 18516 17436
rect 18452 17376 18516 17380
rect 1552 16892 1616 16896
rect 1552 16836 1556 16892
rect 1556 16836 1612 16892
rect 1612 16836 1616 16892
rect 1552 16832 1616 16836
rect 1632 16892 1696 16896
rect 1632 16836 1636 16892
rect 1636 16836 1692 16892
rect 1692 16836 1696 16892
rect 1632 16832 1696 16836
rect 1712 16892 1776 16896
rect 1712 16836 1716 16892
rect 1716 16836 1772 16892
rect 1772 16836 1776 16892
rect 1712 16832 1776 16836
rect 1792 16892 1856 16896
rect 1792 16836 1796 16892
rect 1796 16836 1852 16892
rect 1852 16836 1856 16892
rect 1792 16832 1856 16836
rect 5552 16892 5616 16896
rect 5552 16836 5556 16892
rect 5556 16836 5612 16892
rect 5612 16836 5616 16892
rect 5552 16832 5616 16836
rect 5632 16892 5696 16896
rect 5632 16836 5636 16892
rect 5636 16836 5692 16892
rect 5692 16836 5696 16892
rect 5632 16832 5696 16836
rect 5712 16892 5776 16896
rect 5712 16836 5716 16892
rect 5716 16836 5772 16892
rect 5772 16836 5776 16892
rect 5712 16832 5776 16836
rect 5792 16892 5856 16896
rect 5792 16836 5796 16892
rect 5796 16836 5852 16892
rect 5852 16836 5856 16892
rect 5792 16832 5856 16836
rect 9552 16892 9616 16896
rect 9552 16836 9556 16892
rect 9556 16836 9612 16892
rect 9612 16836 9616 16892
rect 9552 16832 9616 16836
rect 9632 16892 9696 16896
rect 9632 16836 9636 16892
rect 9636 16836 9692 16892
rect 9692 16836 9696 16892
rect 9632 16832 9696 16836
rect 9712 16892 9776 16896
rect 9712 16836 9716 16892
rect 9716 16836 9772 16892
rect 9772 16836 9776 16892
rect 9712 16832 9776 16836
rect 9792 16892 9856 16896
rect 9792 16836 9796 16892
rect 9796 16836 9852 16892
rect 9852 16836 9856 16892
rect 9792 16832 9856 16836
rect 13552 16892 13616 16896
rect 13552 16836 13556 16892
rect 13556 16836 13612 16892
rect 13612 16836 13616 16892
rect 13552 16832 13616 16836
rect 13632 16892 13696 16896
rect 13632 16836 13636 16892
rect 13636 16836 13692 16892
rect 13692 16836 13696 16892
rect 13632 16832 13696 16836
rect 13712 16892 13776 16896
rect 13712 16836 13716 16892
rect 13716 16836 13772 16892
rect 13772 16836 13776 16892
rect 13712 16832 13776 16836
rect 13792 16892 13856 16896
rect 13792 16836 13796 16892
rect 13796 16836 13852 16892
rect 13852 16836 13856 16892
rect 13792 16832 13856 16836
rect 17552 16892 17616 16896
rect 17552 16836 17556 16892
rect 17556 16836 17612 16892
rect 17612 16836 17616 16892
rect 17552 16832 17616 16836
rect 17632 16892 17696 16896
rect 17632 16836 17636 16892
rect 17636 16836 17692 16892
rect 17692 16836 17696 16892
rect 17632 16832 17696 16836
rect 17712 16892 17776 16896
rect 17712 16836 17716 16892
rect 17716 16836 17772 16892
rect 17772 16836 17776 16892
rect 17712 16832 17776 16836
rect 17792 16892 17856 16896
rect 17792 16836 17796 16892
rect 17796 16836 17852 16892
rect 17852 16836 17856 16892
rect 17792 16832 17856 16836
rect 2212 16348 2276 16352
rect 2212 16292 2216 16348
rect 2216 16292 2272 16348
rect 2272 16292 2276 16348
rect 2212 16288 2276 16292
rect 2292 16348 2356 16352
rect 2292 16292 2296 16348
rect 2296 16292 2352 16348
rect 2352 16292 2356 16348
rect 2292 16288 2356 16292
rect 2372 16348 2436 16352
rect 2372 16292 2376 16348
rect 2376 16292 2432 16348
rect 2432 16292 2436 16348
rect 2372 16288 2436 16292
rect 2452 16348 2516 16352
rect 2452 16292 2456 16348
rect 2456 16292 2512 16348
rect 2512 16292 2516 16348
rect 2452 16288 2516 16292
rect 6212 16348 6276 16352
rect 6212 16292 6216 16348
rect 6216 16292 6272 16348
rect 6272 16292 6276 16348
rect 6212 16288 6276 16292
rect 6292 16348 6356 16352
rect 6292 16292 6296 16348
rect 6296 16292 6352 16348
rect 6352 16292 6356 16348
rect 6292 16288 6356 16292
rect 6372 16348 6436 16352
rect 6372 16292 6376 16348
rect 6376 16292 6432 16348
rect 6432 16292 6436 16348
rect 6372 16288 6436 16292
rect 6452 16348 6516 16352
rect 6452 16292 6456 16348
rect 6456 16292 6512 16348
rect 6512 16292 6516 16348
rect 6452 16288 6516 16292
rect 10212 16348 10276 16352
rect 10212 16292 10216 16348
rect 10216 16292 10272 16348
rect 10272 16292 10276 16348
rect 10212 16288 10276 16292
rect 10292 16348 10356 16352
rect 10292 16292 10296 16348
rect 10296 16292 10352 16348
rect 10352 16292 10356 16348
rect 10292 16288 10356 16292
rect 10372 16348 10436 16352
rect 10372 16292 10376 16348
rect 10376 16292 10432 16348
rect 10432 16292 10436 16348
rect 10372 16288 10436 16292
rect 10452 16348 10516 16352
rect 10452 16292 10456 16348
rect 10456 16292 10512 16348
rect 10512 16292 10516 16348
rect 10452 16288 10516 16292
rect 14212 16348 14276 16352
rect 14212 16292 14216 16348
rect 14216 16292 14272 16348
rect 14272 16292 14276 16348
rect 14212 16288 14276 16292
rect 14292 16348 14356 16352
rect 14292 16292 14296 16348
rect 14296 16292 14352 16348
rect 14352 16292 14356 16348
rect 14292 16288 14356 16292
rect 14372 16348 14436 16352
rect 14372 16292 14376 16348
rect 14376 16292 14432 16348
rect 14432 16292 14436 16348
rect 14372 16288 14436 16292
rect 14452 16348 14516 16352
rect 14452 16292 14456 16348
rect 14456 16292 14512 16348
rect 14512 16292 14516 16348
rect 14452 16288 14516 16292
rect 18212 16348 18276 16352
rect 18212 16292 18216 16348
rect 18216 16292 18272 16348
rect 18272 16292 18276 16348
rect 18212 16288 18276 16292
rect 18292 16348 18356 16352
rect 18292 16292 18296 16348
rect 18296 16292 18352 16348
rect 18352 16292 18356 16348
rect 18292 16288 18356 16292
rect 18372 16348 18436 16352
rect 18372 16292 18376 16348
rect 18376 16292 18432 16348
rect 18432 16292 18436 16348
rect 18372 16288 18436 16292
rect 18452 16348 18516 16352
rect 18452 16292 18456 16348
rect 18456 16292 18512 16348
rect 18512 16292 18516 16348
rect 18452 16288 18516 16292
rect 1552 15804 1616 15808
rect 1552 15748 1556 15804
rect 1556 15748 1612 15804
rect 1612 15748 1616 15804
rect 1552 15744 1616 15748
rect 1632 15804 1696 15808
rect 1632 15748 1636 15804
rect 1636 15748 1692 15804
rect 1692 15748 1696 15804
rect 1632 15744 1696 15748
rect 1712 15804 1776 15808
rect 1712 15748 1716 15804
rect 1716 15748 1772 15804
rect 1772 15748 1776 15804
rect 1712 15744 1776 15748
rect 1792 15804 1856 15808
rect 1792 15748 1796 15804
rect 1796 15748 1852 15804
rect 1852 15748 1856 15804
rect 1792 15744 1856 15748
rect 5552 15804 5616 15808
rect 5552 15748 5556 15804
rect 5556 15748 5612 15804
rect 5612 15748 5616 15804
rect 5552 15744 5616 15748
rect 5632 15804 5696 15808
rect 5632 15748 5636 15804
rect 5636 15748 5692 15804
rect 5692 15748 5696 15804
rect 5632 15744 5696 15748
rect 5712 15804 5776 15808
rect 5712 15748 5716 15804
rect 5716 15748 5772 15804
rect 5772 15748 5776 15804
rect 5712 15744 5776 15748
rect 5792 15804 5856 15808
rect 5792 15748 5796 15804
rect 5796 15748 5852 15804
rect 5852 15748 5856 15804
rect 5792 15744 5856 15748
rect 9552 15804 9616 15808
rect 9552 15748 9556 15804
rect 9556 15748 9612 15804
rect 9612 15748 9616 15804
rect 9552 15744 9616 15748
rect 9632 15804 9696 15808
rect 9632 15748 9636 15804
rect 9636 15748 9692 15804
rect 9692 15748 9696 15804
rect 9632 15744 9696 15748
rect 9712 15804 9776 15808
rect 9712 15748 9716 15804
rect 9716 15748 9772 15804
rect 9772 15748 9776 15804
rect 9712 15744 9776 15748
rect 9792 15804 9856 15808
rect 9792 15748 9796 15804
rect 9796 15748 9852 15804
rect 9852 15748 9856 15804
rect 9792 15744 9856 15748
rect 13552 15804 13616 15808
rect 13552 15748 13556 15804
rect 13556 15748 13612 15804
rect 13612 15748 13616 15804
rect 13552 15744 13616 15748
rect 13632 15804 13696 15808
rect 13632 15748 13636 15804
rect 13636 15748 13692 15804
rect 13692 15748 13696 15804
rect 13632 15744 13696 15748
rect 13712 15804 13776 15808
rect 13712 15748 13716 15804
rect 13716 15748 13772 15804
rect 13772 15748 13776 15804
rect 13712 15744 13776 15748
rect 13792 15804 13856 15808
rect 13792 15748 13796 15804
rect 13796 15748 13852 15804
rect 13852 15748 13856 15804
rect 13792 15744 13856 15748
rect 17552 15804 17616 15808
rect 17552 15748 17556 15804
rect 17556 15748 17612 15804
rect 17612 15748 17616 15804
rect 17552 15744 17616 15748
rect 17632 15804 17696 15808
rect 17632 15748 17636 15804
rect 17636 15748 17692 15804
rect 17692 15748 17696 15804
rect 17632 15744 17696 15748
rect 17712 15804 17776 15808
rect 17712 15748 17716 15804
rect 17716 15748 17772 15804
rect 17772 15748 17776 15804
rect 17712 15744 17776 15748
rect 17792 15804 17856 15808
rect 17792 15748 17796 15804
rect 17796 15748 17852 15804
rect 17852 15748 17856 15804
rect 17792 15744 17856 15748
rect 2212 15260 2276 15264
rect 2212 15204 2216 15260
rect 2216 15204 2272 15260
rect 2272 15204 2276 15260
rect 2212 15200 2276 15204
rect 2292 15260 2356 15264
rect 2292 15204 2296 15260
rect 2296 15204 2352 15260
rect 2352 15204 2356 15260
rect 2292 15200 2356 15204
rect 2372 15260 2436 15264
rect 2372 15204 2376 15260
rect 2376 15204 2432 15260
rect 2432 15204 2436 15260
rect 2372 15200 2436 15204
rect 2452 15260 2516 15264
rect 2452 15204 2456 15260
rect 2456 15204 2512 15260
rect 2512 15204 2516 15260
rect 2452 15200 2516 15204
rect 6212 15260 6276 15264
rect 6212 15204 6216 15260
rect 6216 15204 6272 15260
rect 6272 15204 6276 15260
rect 6212 15200 6276 15204
rect 6292 15260 6356 15264
rect 6292 15204 6296 15260
rect 6296 15204 6352 15260
rect 6352 15204 6356 15260
rect 6292 15200 6356 15204
rect 6372 15260 6436 15264
rect 6372 15204 6376 15260
rect 6376 15204 6432 15260
rect 6432 15204 6436 15260
rect 6372 15200 6436 15204
rect 6452 15260 6516 15264
rect 6452 15204 6456 15260
rect 6456 15204 6512 15260
rect 6512 15204 6516 15260
rect 6452 15200 6516 15204
rect 10212 15260 10276 15264
rect 10212 15204 10216 15260
rect 10216 15204 10272 15260
rect 10272 15204 10276 15260
rect 10212 15200 10276 15204
rect 10292 15260 10356 15264
rect 10292 15204 10296 15260
rect 10296 15204 10352 15260
rect 10352 15204 10356 15260
rect 10292 15200 10356 15204
rect 10372 15260 10436 15264
rect 10372 15204 10376 15260
rect 10376 15204 10432 15260
rect 10432 15204 10436 15260
rect 10372 15200 10436 15204
rect 10452 15260 10516 15264
rect 10452 15204 10456 15260
rect 10456 15204 10512 15260
rect 10512 15204 10516 15260
rect 10452 15200 10516 15204
rect 14212 15260 14276 15264
rect 14212 15204 14216 15260
rect 14216 15204 14272 15260
rect 14272 15204 14276 15260
rect 14212 15200 14276 15204
rect 14292 15260 14356 15264
rect 14292 15204 14296 15260
rect 14296 15204 14352 15260
rect 14352 15204 14356 15260
rect 14292 15200 14356 15204
rect 14372 15260 14436 15264
rect 14372 15204 14376 15260
rect 14376 15204 14432 15260
rect 14432 15204 14436 15260
rect 14372 15200 14436 15204
rect 14452 15260 14516 15264
rect 14452 15204 14456 15260
rect 14456 15204 14512 15260
rect 14512 15204 14516 15260
rect 14452 15200 14516 15204
rect 18212 15260 18276 15264
rect 18212 15204 18216 15260
rect 18216 15204 18272 15260
rect 18272 15204 18276 15260
rect 18212 15200 18276 15204
rect 18292 15260 18356 15264
rect 18292 15204 18296 15260
rect 18296 15204 18352 15260
rect 18352 15204 18356 15260
rect 18292 15200 18356 15204
rect 18372 15260 18436 15264
rect 18372 15204 18376 15260
rect 18376 15204 18432 15260
rect 18432 15204 18436 15260
rect 18372 15200 18436 15204
rect 18452 15260 18516 15264
rect 18452 15204 18456 15260
rect 18456 15204 18512 15260
rect 18512 15204 18516 15260
rect 18452 15200 18516 15204
rect 1552 14716 1616 14720
rect 1552 14660 1556 14716
rect 1556 14660 1612 14716
rect 1612 14660 1616 14716
rect 1552 14656 1616 14660
rect 1632 14716 1696 14720
rect 1632 14660 1636 14716
rect 1636 14660 1692 14716
rect 1692 14660 1696 14716
rect 1632 14656 1696 14660
rect 1712 14716 1776 14720
rect 1712 14660 1716 14716
rect 1716 14660 1772 14716
rect 1772 14660 1776 14716
rect 1712 14656 1776 14660
rect 1792 14716 1856 14720
rect 1792 14660 1796 14716
rect 1796 14660 1852 14716
rect 1852 14660 1856 14716
rect 1792 14656 1856 14660
rect 5552 14716 5616 14720
rect 5552 14660 5556 14716
rect 5556 14660 5612 14716
rect 5612 14660 5616 14716
rect 5552 14656 5616 14660
rect 5632 14716 5696 14720
rect 5632 14660 5636 14716
rect 5636 14660 5692 14716
rect 5692 14660 5696 14716
rect 5632 14656 5696 14660
rect 5712 14716 5776 14720
rect 5712 14660 5716 14716
rect 5716 14660 5772 14716
rect 5772 14660 5776 14716
rect 5712 14656 5776 14660
rect 5792 14716 5856 14720
rect 5792 14660 5796 14716
rect 5796 14660 5852 14716
rect 5852 14660 5856 14716
rect 5792 14656 5856 14660
rect 9552 14716 9616 14720
rect 9552 14660 9556 14716
rect 9556 14660 9612 14716
rect 9612 14660 9616 14716
rect 9552 14656 9616 14660
rect 9632 14716 9696 14720
rect 9632 14660 9636 14716
rect 9636 14660 9692 14716
rect 9692 14660 9696 14716
rect 9632 14656 9696 14660
rect 9712 14716 9776 14720
rect 9712 14660 9716 14716
rect 9716 14660 9772 14716
rect 9772 14660 9776 14716
rect 9712 14656 9776 14660
rect 9792 14716 9856 14720
rect 9792 14660 9796 14716
rect 9796 14660 9852 14716
rect 9852 14660 9856 14716
rect 9792 14656 9856 14660
rect 13552 14716 13616 14720
rect 13552 14660 13556 14716
rect 13556 14660 13612 14716
rect 13612 14660 13616 14716
rect 13552 14656 13616 14660
rect 13632 14716 13696 14720
rect 13632 14660 13636 14716
rect 13636 14660 13692 14716
rect 13692 14660 13696 14716
rect 13632 14656 13696 14660
rect 13712 14716 13776 14720
rect 13712 14660 13716 14716
rect 13716 14660 13772 14716
rect 13772 14660 13776 14716
rect 13712 14656 13776 14660
rect 13792 14716 13856 14720
rect 13792 14660 13796 14716
rect 13796 14660 13852 14716
rect 13852 14660 13856 14716
rect 13792 14656 13856 14660
rect 17552 14716 17616 14720
rect 17552 14660 17556 14716
rect 17556 14660 17612 14716
rect 17612 14660 17616 14716
rect 17552 14656 17616 14660
rect 17632 14716 17696 14720
rect 17632 14660 17636 14716
rect 17636 14660 17692 14716
rect 17692 14660 17696 14716
rect 17632 14656 17696 14660
rect 17712 14716 17776 14720
rect 17712 14660 17716 14716
rect 17716 14660 17772 14716
rect 17772 14660 17776 14716
rect 17712 14656 17776 14660
rect 17792 14716 17856 14720
rect 17792 14660 17796 14716
rect 17796 14660 17852 14716
rect 17852 14660 17856 14716
rect 17792 14656 17856 14660
rect 2212 14172 2276 14176
rect 2212 14116 2216 14172
rect 2216 14116 2272 14172
rect 2272 14116 2276 14172
rect 2212 14112 2276 14116
rect 2292 14172 2356 14176
rect 2292 14116 2296 14172
rect 2296 14116 2352 14172
rect 2352 14116 2356 14172
rect 2292 14112 2356 14116
rect 2372 14172 2436 14176
rect 2372 14116 2376 14172
rect 2376 14116 2432 14172
rect 2432 14116 2436 14172
rect 2372 14112 2436 14116
rect 2452 14172 2516 14176
rect 2452 14116 2456 14172
rect 2456 14116 2512 14172
rect 2512 14116 2516 14172
rect 2452 14112 2516 14116
rect 6212 14172 6276 14176
rect 6212 14116 6216 14172
rect 6216 14116 6272 14172
rect 6272 14116 6276 14172
rect 6212 14112 6276 14116
rect 6292 14172 6356 14176
rect 6292 14116 6296 14172
rect 6296 14116 6352 14172
rect 6352 14116 6356 14172
rect 6292 14112 6356 14116
rect 6372 14172 6436 14176
rect 6372 14116 6376 14172
rect 6376 14116 6432 14172
rect 6432 14116 6436 14172
rect 6372 14112 6436 14116
rect 6452 14172 6516 14176
rect 6452 14116 6456 14172
rect 6456 14116 6512 14172
rect 6512 14116 6516 14172
rect 6452 14112 6516 14116
rect 10212 14172 10276 14176
rect 10212 14116 10216 14172
rect 10216 14116 10272 14172
rect 10272 14116 10276 14172
rect 10212 14112 10276 14116
rect 10292 14172 10356 14176
rect 10292 14116 10296 14172
rect 10296 14116 10352 14172
rect 10352 14116 10356 14172
rect 10292 14112 10356 14116
rect 10372 14172 10436 14176
rect 10372 14116 10376 14172
rect 10376 14116 10432 14172
rect 10432 14116 10436 14172
rect 10372 14112 10436 14116
rect 10452 14172 10516 14176
rect 10452 14116 10456 14172
rect 10456 14116 10512 14172
rect 10512 14116 10516 14172
rect 10452 14112 10516 14116
rect 14212 14172 14276 14176
rect 14212 14116 14216 14172
rect 14216 14116 14272 14172
rect 14272 14116 14276 14172
rect 14212 14112 14276 14116
rect 14292 14172 14356 14176
rect 14292 14116 14296 14172
rect 14296 14116 14352 14172
rect 14352 14116 14356 14172
rect 14292 14112 14356 14116
rect 14372 14172 14436 14176
rect 14372 14116 14376 14172
rect 14376 14116 14432 14172
rect 14432 14116 14436 14172
rect 14372 14112 14436 14116
rect 14452 14172 14516 14176
rect 14452 14116 14456 14172
rect 14456 14116 14512 14172
rect 14512 14116 14516 14172
rect 14452 14112 14516 14116
rect 18212 14172 18276 14176
rect 18212 14116 18216 14172
rect 18216 14116 18272 14172
rect 18272 14116 18276 14172
rect 18212 14112 18276 14116
rect 18292 14172 18356 14176
rect 18292 14116 18296 14172
rect 18296 14116 18352 14172
rect 18352 14116 18356 14172
rect 18292 14112 18356 14116
rect 18372 14172 18436 14176
rect 18372 14116 18376 14172
rect 18376 14116 18432 14172
rect 18432 14116 18436 14172
rect 18372 14112 18436 14116
rect 18452 14172 18516 14176
rect 18452 14116 18456 14172
rect 18456 14116 18512 14172
rect 18512 14116 18516 14172
rect 18452 14112 18516 14116
rect 1552 13628 1616 13632
rect 1552 13572 1556 13628
rect 1556 13572 1612 13628
rect 1612 13572 1616 13628
rect 1552 13568 1616 13572
rect 1632 13628 1696 13632
rect 1632 13572 1636 13628
rect 1636 13572 1692 13628
rect 1692 13572 1696 13628
rect 1632 13568 1696 13572
rect 1712 13628 1776 13632
rect 1712 13572 1716 13628
rect 1716 13572 1772 13628
rect 1772 13572 1776 13628
rect 1712 13568 1776 13572
rect 1792 13628 1856 13632
rect 1792 13572 1796 13628
rect 1796 13572 1852 13628
rect 1852 13572 1856 13628
rect 1792 13568 1856 13572
rect 5552 13628 5616 13632
rect 5552 13572 5556 13628
rect 5556 13572 5612 13628
rect 5612 13572 5616 13628
rect 5552 13568 5616 13572
rect 5632 13628 5696 13632
rect 5632 13572 5636 13628
rect 5636 13572 5692 13628
rect 5692 13572 5696 13628
rect 5632 13568 5696 13572
rect 5712 13628 5776 13632
rect 5712 13572 5716 13628
rect 5716 13572 5772 13628
rect 5772 13572 5776 13628
rect 5712 13568 5776 13572
rect 5792 13628 5856 13632
rect 5792 13572 5796 13628
rect 5796 13572 5852 13628
rect 5852 13572 5856 13628
rect 5792 13568 5856 13572
rect 9552 13628 9616 13632
rect 9552 13572 9556 13628
rect 9556 13572 9612 13628
rect 9612 13572 9616 13628
rect 9552 13568 9616 13572
rect 9632 13628 9696 13632
rect 9632 13572 9636 13628
rect 9636 13572 9692 13628
rect 9692 13572 9696 13628
rect 9632 13568 9696 13572
rect 9712 13628 9776 13632
rect 9712 13572 9716 13628
rect 9716 13572 9772 13628
rect 9772 13572 9776 13628
rect 9712 13568 9776 13572
rect 9792 13628 9856 13632
rect 9792 13572 9796 13628
rect 9796 13572 9852 13628
rect 9852 13572 9856 13628
rect 9792 13568 9856 13572
rect 13552 13628 13616 13632
rect 13552 13572 13556 13628
rect 13556 13572 13612 13628
rect 13612 13572 13616 13628
rect 13552 13568 13616 13572
rect 13632 13628 13696 13632
rect 13632 13572 13636 13628
rect 13636 13572 13692 13628
rect 13692 13572 13696 13628
rect 13632 13568 13696 13572
rect 13712 13628 13776 13632
rect 13712 13572 13716 13628
rect 13716 13572 13772 13628
rect 13772 13572 13776 13628
rect 13712 13568 13776 13572
rect 13792 13628 13856 13632
rect 13792 13572 13796 13628
rect 13796 13572 13852 13628
rect 13852 13572 13856 13628
rect 13792 13568 13856 13572
rect 17552 13628 17616 13632
rect 17552 13572 17556 13628
rect 17556 13572 17612 13628
rect 17612 13572 17616 13628
rect 17552 13568 17616 13572
rect 17632 13628 17696 13632
rect 17632 13572 17636 13628
rect 17636 13572 17692 13628
rect 17692 13572 17696 13628
rect 17632 13568 17696 13572
rect 17712 13628 17776 13632
rect 17712 13572 17716 13628
rect 17716 13572 17772 13628
rect 17772 13572 17776 13628
rect 17712 13568 17776 13572
rect 17792 13628 17856 13632
rect 17792 13572 17796 13628
rect 17796 13572 17852 13628
rect 17852 13572 17856 13628
rect 17792 13568 17856 13572
rect 2212 13084 2276 13088
rect 2212 13028 2216 13084
rect 2216 13028 2272 13084
rect 2272 13028 2276 13084
rect 2212 13024 2276 13028
rect 2292 13084 2356 13088
rect 2292 13028 2296 13084
rect 2296 13028 2352 13084
rect 2352 13028 2356 13084
rect 2292 13024 2356 13028
rect 2372 13084 2436 13088
rect 2372 13028 2376 13084
rect 2376 13028 2432 13084
rect 2432 13028 2436 13084
rect 2372 13024 2436 13028
rect 2452 13084 2516 13088
rect 2452 13028 2456 13084
rect 2456 13028 2512 13084
rect 2512 13028 2516 13084
rect 2452 13024 2516 13028
rect 6212 13084 6276 13088
rect 6212 13028 6216 13084
rect 6216 13028 6272 13084
rect 6272 13028 6276 13084
rect 6212 13024 6276 13028
rect 6292 13084 6356 13088
rect 6292 13028 6296 13084
rect 6296 13028 6352 13084
rect 6352 13028 6356 13084
rect 6292 13024 6356 13028
rect 6372 13084 6436 13088
rect 6372 13028 6376 13084
rect 6376 13028 6432 13084
rect 6432 13028 6436 13084
rect 6372 13024 6436 13028
rect 6452 13084 6516 13088
rect 6452 13028 6456 13084
rect 6456 13028 6512 13084
rect 6512 13028 6516 13084
rect 6452 13024 6516 13028
rect 10212 13084 10276 13088
rect 10212 13028 10216 13084
rect 10216 13028 10272 13084
rect 10272 13028 10276 13084
rect 10212 13024 10276 13028
rect 10292 13084 10356 13088
rect 10292 13028 10296 13084
rect 10296 13028 10352 13084
rect 10352 13028 10356 13084
rect 10292 13024 10356 13028
rect 10372 13084 10436 13088
rect 10372 13028 10376 13084
rect 10376 13028 10432 13084
rect 10432 13028 10436 13084
rect 10372 13024 10436 13028
rect 10452 13084 10516 13088
rect 10452 13028 10456 13084
rect 10456 13028 10512 13084
rect 10512 13028 10516 13084
rect 10452 13024 10516 13028
rect 14212 13084 14276 13088
rect 14212 13028 14216 13084
rect 14216 13028 14272 13084
rect 14272 13028 14276 13084
rect 14212 13024 14276 13028
rect 14292 13084 14356 13088
rect 14292 13028 14296 13084
rect 14296 13028 14352 13084
rect 14352 13028 14356 13084
rect 14292 13024 14356 13028
rect 14372 13084 14436 13088
rect 14372 13028 14376 13084
rect 14376 13028 14432 13084
rect 14432 13028 14436 13084
rect 14372 13024 14436 13028
rect 14452 13084 14516 13088
rect 14452 13028 14456 13084
rect 14456 13028 14512 13084
rect 14512 13028 14516 13084
rect 14452 13024 14516 13028
rect 18212 13084 18276 13088
rect 18212 13028 18216 13084
rect 18216 13028 18272 13084
rect 18272 13028 18276 13084
rect 18212 13024 18276 13028
rect 18292 13084 18356 13088
rect 18292 13028 18296 13084
rect 18296 13028 18352 13084
rect 18352 13028 18356 13084
rect 18292 13024 18356 13028
rect 18372 13084 18436 13088
rect 18372 13028 18376 13084
rect 18376 13028 18432 13084
rect 18432 13028 18436 13084
rect 18372 13024 18436 13028
rect 18452 13084 18516 13088
rect 18452 13028 18456 13084
rect 18456 13028 18512 13084
rect 18512 13028 18516 13084
rect 18452 13024 18516 13028
rect 1552 12540 1616 12544
rect 1552 12484 1556 12540
rect 1556 12484 1612 12540
rect 1612 12484 1616 12540
rect 1552 12480 1616 12484
rect 1632 12540 1696 12544
rect 1632 12484 1636 12540
rect 1636 12484 1692 12540
rect 1692 12484 1696 12540
rect 1632 12480 1696 12484
rect 1712 12540 1776 12544
rect 1712 12484 1716 12540
rect 1716 12484 1772 12540
rect 1772 12484 1776 12540
rect 1712 12480 1776 12484
rect 1792 12540 1856 12544
rect 1792 12484 1796 12540
rect 1796 12484 1852 12540
rect 1852 12484 1856 12540
rect 1792 12480 1856 12484
rect 5552 12540 5616 12544
rect 5552 12484 5556 12540
rect 5556 12484 5612 12540
rect 5612 12484 5616 12540
rect 5552 12480 5616 12484
rect 5632 12540 5696 12544
rect 5632 12484 5636 12540
rect 5636 12484 5692 12540
rect 5692 12484 5696 12540
rect 5632 12480 5696 12484
rect 5712 12540 5776 12544
rect 5712 12484 5716 12540
rect 5716 12484 5772 12540
rect 5772 12484 5776 12540
rect 5712 12480 5776 12484
rect 5792 12540 5856 12544
rect 5792 12484 5796 12540
rect 5796 12484 5852 12540
rect 5852 12484 5856 12540
rect 5792 12480 5856 12484
rect 9552 12540 9616 12544
rect 9552 12484 9556 12540
rect 9556 12484 9612 12540
rect 9612 12484 9616 12540
rect 9552 12480 9616 12484
rect 9632 12540 9696 12544
rect 9632 12484 9636 12540
rect 9636 12484 9692 12540
rect 9692 12484 9696 12540
rect 9632 12480 9696 12484
rect 9712 12540 9776 12544
rect 9712 12484 9716 12540
rect 9716 12484 9772 12540
rect 9772 12484 9776 12540
rect 9712 12480 9776 12484
rect 9792 12540 9856 12544
rect 9792 12484 9796 12540
rect 9796 12484 9852 12540
rect 9852 12484 9856 12540
rect 9792 12480 9856 12484
rect 13552 12540 13616 12544
rect 13552 12484 13556 12540
rect 13556 12484 13612 12540
rect 13612 12484 13616 12540
rect 13552 12480 13616 12484
rect 13632 12540 13696 12544
rect 13632 12484 13636 12540
rect 13636 12484 13692 12540
rect 13692 12484 13696 12540
rect 13632 12480 13696 12484
rect 13712 12540 13776 12544
rect 13712 12484 13716 12540
rect 13716 12484 13772 12540
rect 13772 12484 13776 12540
rect 13712 12480 13776 12484
rect 13792 12540 13856 12544
rect 13792 12484 13796 12540
rect 13796 12484 13852 12540
rect 13852 12484 13856 12540
rect 13792 12480 13856 12484
rect 17552 12540 17616 12544
rect 17552 12484 17556 12540
rect 17556 12484 17612 12540
rect 17612 12484 17616 12540
rect 17552 12480 17616 12484
rect 17632 12540 17696 12544
rect 17632 12484 17636 12540
rect 17636 12484 17692 12540
rect 17692 12484 17696 12540
rect 17632 12480 17696 12484
rect 17712 12540 17776 12544
rect 17712 12484 17716 12540
rect 17716 12484 17772 12540
rect 17772 12484 17776 12540
rect 17712 12480 17776 12484
rect 17792 12540 17856 12544
rect 17792 12484 17796 12540
rect 17796 12484 17852 12540
rect 17852 12484 17856 12540
rect 17792 12480 17856 12484
rect 2212 11996 2276 12000
rect 2212 11940 2216 11996
rect 2216 11940 2272 11996
rect 2272 11940 2276 11996
rect 2212 11936 2276 11940
rect 2292 11996 2356 12000
rect 2292 11940 2296 11996
rect 2296 11940 2352 11996
rect 2352 11940 2356 11996
rect 2292 11936 2356 11940
rect 2372 11996 2436 12000
rect 2372 11940 2376 11996
rect 2376 11940 2432 11996
rect 2432 11940 2436 11996
rect 2372 11936 2436 11940
rect 2452 11996 2516 12000
rect 2452 11940 2456 11996
rect 2456 11940 2512 11996
rect 2512 11940 2516 11996
rect 2452 11936 2516 11940
rect 6212 11996 6276 12000
rect 6212 11940 6216 11996
rect 6216 11940 6272 11996
rect 6272 11940 6276 11996
rect 6212 11936 6276 11940
rect 6292 11996 6356 12000
rect 6292 11940 6296 11996
rect 6296 11940 6352 11996
rect 6352 11940 6356 11996
rect 6292 11936 6356 11940
rect 6372 11996 6436 12000
rect 6372 11940 6376 11996
rect 6376 11940 6432 11996
rect 6432 11940 6436 11996
rect 6372 11936 6436 11940
rect 6452 11996 6516 12000
rect 6452 11940 6456 11996
rect 6456 11940 6512 11996
rect 6512 11940 6516 11996
rect 6452 11936 6516 11940
rect 10212 11996 10276 12000
rect 10212 11940 10216 11996
rect 10216 11940 10272 11996
rect 10272 11940 10276 11996
rect 10212 11936 10276 11940
rect 10292 11996 10356 12000
rect 10292 11940 10296 11996
rect 10296 11940 10352 11996
rect 10352 11940 10356 11996
rect 10292 11936 10356 11940
rect 10372 11996 10436 12000
rect 10372 11940 10376 11996
rect 10376 11940 10432 11996
rect 10432 11940 10436 11996
rect 10372 11936 10436 11940
rect 10452 11996 10516 12000
rect 10452 11940 10456 11996
rect 10456 11940 10512 11996
rect 10512 11940 10516 11996
rect 10452 11936 10516 11940
rect 14212 11996 14276 12000
rect 14212 11940 14216 11996
rect 14216 11940 14272 11996
rect 14272 11940 14276 11996
rect 14212 11936 14276 11940
rect 14292 11996 14356 12000
rect 14292 11940 14296 11996
rect 14296 11940 14352 11996
rect 14352 11940 14356 11996
rect 14292 11936 14356 11940
rect 14372 11996 14436 12000
rect 14372 11940 14376 11996
rect 14376 11940 14432 11996
rect 14432 11940 14436 11996
rect 14372 11936 14436 11940
rect 14452 11996 14516 12000
rect 14452 11940 14456 11996
rect 14456 11940 14512 11996
rect 14512 11940 14516 11996
rect 14452 11936 14516 11940
rect 18212 11996 18276 12000
rect 18212 11940 18216 11996
rect 18216 11940 18272 11996
rect 18272 11940 18276 11996
rect 18212 11936 18276 11940
rect 18292 11996 18356 12000
rect 18292 11940 18296 11996
rect 18296 11940 18352 11996
rect 18352 11940 18356 11996
rect 18292 11936 18356 11940
rect 18372 11996 18436 12000
rect 18372 11940 18376 11996
rect 18376 11940 18432 11996
rect 18432 11940 18436 11996
rect 18372 11936 18436 11940
rect 18452 11996 18516 12000
rect 18452 11940 18456 11996
rect 18456 11940 18512 11996
rect 18512 11940 18516 11996
rect 18452 11936 18516 11940
rect 1552 11452 1616 11456
rect 1552 11396 1556 11452
rect 1556 11396 1612 11452
rect 1612 11396 1616 11452
rect 1552 11392 1616 11396
rect 1632 11452 1696 11456
rect 1632 11396 1636 11452
rect 1636 11396 1692 11452
rect 1692 11396 1696 11452
rect 1632 11392 1696 11396
rect 1712 11452 1776 11456
rect 1712 11396 1716 11452
rect 1716 11396 1772 11452
rect 1772 11396 1776 11452
rect 1712 11392 1776 11396
rect 1792 11452 1856 11456
rect 1792 11396 1796 11452
rect 1796 11396 1852 11452
rect 1852 11396 1856 11452
rect 1792 11392 1856 11396
rect 5552 11452 5616 11456
rect 5552 11396 5556 11452
rect 5556 11396 5612 11452
rect 5612 11396 5616 11452
rect 5552 11392 5616 11396
rect 5632 11452 5696 11456
rect 5632 11396 5636 11452
rect 5636 11396 5692 11452
rect 5692 11396 5696 11452
rect 5632 11392 5696 11396
rect 5712 11452 5776 11456
rect 5712 11396 5716 11452
rect 5716 11396 5772 11452
rect 5772 11396 5776 11452
rect 5712 11392 5776 11396
rect 5792 11452 5856 11456
rect 5792 11396 5796 11452
rect 5796 11396 5852 11452
rect 5852 11396 5856 11452
rect 5792 11392 5856 11396
rect 9552 11452 9616 11456
rect 9552 11396 9556 11452
rect 9556 11396 9612 11452
rect 9612 11396 9616 11452
rect 9552 11392 9616 11396
rect 9632 11452 9696 11456
rect 9632 11396 9636 11452
rect 9636 11396 9692 11452
rect 9692 11396 9696 11452
rect 9632 11392 9696 11396
rect 9712 11452 9776 11456
rect 9712 11396 9716 11452
rect 9716 11396 9772 11452
rect 9772 11396 9776 11452
rect 9712 11392 9776 11396
rect 9792 11452 9856 11456
rect 9792 11396 9796 11452
rect 9796 11396 9852 11452
rect 9852 11396 9856 11452
rect 9792 11392 9856 11396
rect 13552 11452 13616 11456
rect 13552 11396 13556 11452
rect 13556 11396 13612 11452
rect 13612 11396 13616 11452
rect 13552 11392 13616 11396
rect 13632 11452 13696 11456
rect 13632 11396 13636 11452
rect 13636 11396 13692 11452
rect 13692 11396 13696 11452
rect 13632 11392 13696 11396
rect 13712 11452 13776 11456
rect 13712 11396 13716 11452
rect 13716 11396 13772 11452
rect 13772 11396 13776 11452
rect 13712 11392 13776 11396
rect 13792 11452 13856 11456
rect 13792 11396 13796 11452
rect 13796 11396 13852 11452
rect 13852 11396 13856 11452
rect 13792 11392 13856 11396
rect 17552 11452 17616 11456
rect 17552 11396 17556 11452
rect 17556 11396 17612 11452
rect 17612 11396 17616 11452
rect 17552 11392 17616 11396
rect 17632 11452 17696 11456
rect 17632 11396 17636 11452
rect 17636 11396 17692 11452
rect 17692 11396 17696 11452
rect 17632 11392 17696 11396
rect 17712 11452 17776 11456
rect 17712 11396 17716 11452
rect 17716 11396 17772 11452
rect 17772 11396 17776 11452
rect 17712 11392 17776 11396
rect 17792 11452 17856 11456
rect 17792 11396 17796 11452
rect 17796 11396 17852 11452
rect 17852 11396 17856 11452
rect 17792 11392 17856 11396
rect 2212 10908 2276 10912
rect 2212 10852 2216 10908
rect 2216 10852 2272 10908
rect 2272 10852 2276 10908
rect 2212 10848 2276 10852
rect 2292 10908 2356 10912
rect 2292 10852 2296 10908
rect 2296 10852 2352 10908
rect 2352 10852 2356 10908
rect 2292 10848 2356 10852
rect 2372 10908 2436 10912
rect 2372 10852 2376 10908
rect 2376 10852 2432 10908
rect 2432 10852 2436 10908
rect 2372 10848 2436 10852
rect 2452 10908 2516 10912
rect 2452 10852 2456 10908
rect 2456 10852 2512 10908
rect 2512 10852 2516 10908
rect 2452 10848 2516 10852
rect 6212 10908 6276 10912
rect 6212 10852 6216 10908
rect 6216 10852 6272 10908
rect 6272 10852 6276 10908
rect 6212 10848 6276 10852
rect 6292 10908 6356 10912
rect 6292 10852 6296 10908
rect 6296 10852 6352 10908
rect 6352 10852 6356 10908
rect 6292 10848 6356 10852
rect 6372 10908 6436 10912
rect 6372 10852 6376 10908
rect 6376 10852 6432 10908
rect 6432 10852 6436 10908
rect 6372 10848 6436 10852
rect 6452 10908 6516 10912
rect 6452 10852 6456 10908
rect 6456 10852 6512 10908
rect 6512 10852 6516 10908
rect 6452 10848 6516 10852
rect 10212 10908 10276 10912
rect 10212 10852 10216 10908
rect 10216 10852 10272 10908
rect 10272 10852 10276 10908
rect 10212 10848 10276 10852
rect 10292 10908 10356 10912
rect 10292 10852 10296 10908
rect 10296 10852 10352 10908
rect 10352 10852 10356 10908
rect 10292 10848 10356 10852
rect 10372 10908 10436 10912
rect 10372 10852 10376 10908
rect 10376 10852 10432 10908
rect 10432 10852 10436 10908
rect 10372 10848 10436 10852
rect 10452 10908 10516 10912
rect 10452 10852 10456 10908
rect 10456 10852 10512 10908
rect 10512 10852 10516 10908
rect 10452 10848 10516 10852
rect 14212 10908 14276 10912
rect 14212 10852 14216 10908
rect 14216 10852 14272 10908
rect 14272 10852 14276 10908
rect 14212 10848 14276 10852
rect 14292 10908 14356 10912
rect 14292 10852 14296 10908
rect 14296 10852 14352 10908
rect 14352 10852 14356 10908
rect 14292 10848 14356 10852
rect 14372 10908 14436 10912
rect 14372 10852 14376 10908
rect 14376 10852 14432 10908
rect 14432 10852 14436 10908
rect 14372 10848 14436 10852
rect 14452 10908 14516 10912
rect 14452 10852 14456 10908
rect 14456 10852 14512 10908
rect 14512 10852 14516 10908
rect 14452 10848 14516 10852
rect 18212 10908 18276 10912
rect 18212 10852 18216 10908
rect 18216 10852 18272 10908
rect 18272 10852 18276 10908
rect 18212 10848 18276 10852
rect 18292 10908 18356 10912
rect 18292 10852 18296 10908
rect 18296 10852 18352 10908
rect 18352 10852 18356 10908
rect 18292 10848 18356 10852
rect 18372 10908 18436 10912
rect 18372 10852 18376 10908
rect 18376 10852 18432 10908
rect 18432 10852 18436 10908
rect 18372 10848 18436 10852
rect 18452 10908 18516 10912
rect 18452 10852 18456 10908
rect 18456 10852 18512 10908
rect 18512 10852 18516 10908
rect 18452 10848 18516 10852
rect 1552 10364 1616 10368
rect 1552 10308 1556 10364
rect 1556 10308 1612 10364
rect 1612 10308 1616 10364
rect 1552 10304 1616 10308
rect 1632 10364 1696 10368
rect 1632 10308 1636 10364
rect 1636 10308 1692 10364
rect 1692 10308 1696 10364
rect 1632 10304 1696 10308
rect 1712 10364 1776 10368
rect 1712 10308 1716 10364
rect 1716 10308 1772 10364
rect 1772 10308 1776 10364
rect 1712 10304 1776 10308
rect 1792 10364 1856 10368
rect 1792 10308 1796 10364
rect 1796 10308 1852 10364
rect 1852 10308 1856 10364
rect 1792 10304 1856 10308
rect 5552 10364 5616 10368
rect 5552 10308 5556 10364
rect 5556 10308 5612 10364
rect 5612 10308 5616 10364
rect 5552 10304 5616 10308
rect 5632 10364 5696 10368
rect 5632 10308 5636 10364
rect 5636 10308 5692 10364
rect 5692 10308 5696 10364
rect 5632 10304 5696 10308
rect 5712 10364 5776 10368
rect 5712 10308 5716 10364
rect 5716 10308 5772 10364
rect 5772 10308 5776 10364
rect 5712 10304 5776 10308
rect 5792 10364 5856 10368
rect 5792 10308 5796 10364
rect 5796 10308 5852 10364
rect 5852 10308 5856 10364
rect 5792 10304 5856 10308
rect 9552 10364 9616 10368
rect 9552 10308 9556 10364
rect 9556 10308 9612 10364
rect 9612 10308 9616 10364
rect 9552 10304 9616 10308
rect 9632 10364 9696 10368
rect 9632 10308 9636 10364
rect 9636 10308 9692 10364
rect 9692 10308 9696 10364
rect 9632 10304 9696 10308
rect 9712 10364 9776 10368
rect 9712 10308 9716 10364
rect 9716 10308 9772 10364
rect 9772 10308 9776 10364
rect 9712 10304 9776 10308
rect 9792 10364 9856 10368
rect 9792 10308 9796 10364
rect 9796 10308 9852 10364
rect 9852 10308 9856 10364
rect 9792 10304 9856 10308
rect 13552 10364 13616 10368
rect 13552 10308 13556 10364
rect 13556 10308 13612 10364
rect 13612 10308 13616 10364
rect 13552 10304 13616 10308
rect 13632 10364 13696 10368
rect 13632 10308 13636 10364
rect 13636 10308 13692 10364
rect 13692 10308 13696 10364
rect 13632 10304 13696 10308
rect 13712 10364 13776 10368
rect 13712 10308 13716 10364
rect 13716 10308 13772 10364
rect 13772 10308 13776 10364
rect 13712 10304 13776 10308
rect 13792 10364 13856 10368
rect 13792 10308 13796 10364
rect 13796 10308 13852 10364
rect 13852 10308 13856 10364
rect 13792 10304 13856 10308
rect 17552 10364 17616 10368
rect 17552 10308 17556 10364
rect 17556 10308 17612 10364
rect 17612 10308 17616 10364
rect 17552 10304 17616 10308
rect 17632 10364 17696 10368
rect 17632 10308 17636 10364
rect 17636 10308 17692 10364
rect 17692 10308 17696 10364
rect 17632 10304 17696 10308
rect 17712 10364 17776 10368
rect 17712 10308 17716 10364
rect 17716 10308 17772 10364
rect 17772 10308 17776 10364
rect 17712 10304 17776 10308
rect 17792 10364 17856 10368
rect 17792 10308 17796 10364
rect 17796 10308 17852 10364
rect 17852 10308 17856 10364
rect 17792 10304 17856 10308
rect 2212 9820 2276 9824
rect 2212 9764 2216 9820
rect 2216 9764 2272 9820
rect 2272 9764 2276 9820
rect 2212 9760 2276 9764
rect 2292 9820 2356 9824
rect 2292 9764 2296 9820
rect 2296 9764 2352 9820
rect 2352 9764 2356 9820
rect 2292 9760 2356 9764
rect 2372 9820 2436 9824
rect 2372 9764 2376 9820
rect 2376 9764 2432 9820
rect 2432 9764 2436 9820
rect 2372 9760 2436 9764
rect 2452 9820 2516 9824
rect 2452 9764 2456 9820
rect 2456 9764 2512 9820
rect 2512 9764 2516 9820
rect 2452 9760 2516 9764
rect 6212 9820 6276 9824
rect 6212 9764 6216 9820
rect 6216 9764 6272 9820
rect 6272 9764 6276 9820
rect 6212 9760 6276 9764
rect 6292 9820 6356 9824
rect 6292 9764 6296 9820
rect 6296 9764 6352 9820
rect 6352 9764 6356 9820
rect 6292 9760 6356 9764
rect 6372 9820 6436 9824
rect 6372 9764 6376 9820
rect 6376 9764 6432 9820
rect 6432 9764 6436 9820
rect 6372 9760 6436 9764
rect 6452 9820 6516 9824
rect 6452 9764 6456 9820
rect 6456 9764 6512 9820
rect 6512 9764 6516 9820
rect 6452 9760 6516 9764
rect 10212 9820 10276 9824
rect 10212 9764 10216 9820
rect 10216 9764 10272 9820
rect 10272 9764 10276 9820
rect 10212 9760 10276 9764
rect 10292 9820 10356 9824
rect 10292 9764 10296 9820
rect 10296 9764 10352 9820
rect 10352 9764 10356 9820
rect 10292 9760 10356 9764
rect 10372 9820 10436 9824
rect 10372 9764 10376 9820
rect 10376 9764 10432 9820
rect 10432 9764 10436 9820
rect 10372 9760 10436 9764
rect 10452 9820 10516 9824
rect 10452 9764 10456 9820
rect 10456 9764 10512 9820
rect 10512 9764 10516 9820
rect 10452 9760 10516 9764
rect 14212 9820 14276 9824
rect 14212 9764 14216 9820
rect 14216 9764 14272 9820
rect 14272 9764 14276 9820
rect 14212 9760 14276 9764
rect 14292 9820 14356 9824
rect 14292 9764 14296 9820
rect 14296 9764 14352 9820
rect 14352 9764 14356 9820
rect 14292 9760 14356 9764
rect 14372 9820 14436 9824
rect 14372 9764 14376 9820
rect 14376 9764 14432 9820
rect 14432 9764 14436 9820
rect 14372 9760 14436 9764
rect 14452 9820 14516 9824
rect 14452 9764 14456 9820
rect 14456 9764 14512 9820
rect 14512 9764 14516 9820
rect 14452 9760 14516 9764
rect 18212 9820 18276 9824
rect 18212 9764 18216 9820
rect 18216 9764 18272 9820
rect 18272 9764 18276 9820
rect 18212 9760 18276 9764
rect 18292 9820 18356 9824
rect 18292 9764 18296 9820
rect 18296 9764 18352 9820
rect 18352 9764 18356 9820
rect 18292 9760 18356 9764
rect 18372 9820 18436 9824
rect 18372 9764 18376 9820
rect 18376 9764 18432 9820
rect 18432 9764 18436 9820
rect 18372 9760 18436 9764
rect 18452 9820 18516 9824
rect 18452 9764 18456 9820
rect 18456 9764 18512 9820
rect 18512 9764 18516 9820
rect 18452 9760 18516 9764
rect 1552 9276 1616 9280
rect 1552 9220 1556 9276
rect 1556 9220 1612 9276
rect 1612 9220 1616 9276
rect 1552 9216 1616 9220
rect 1632 9276 1696 9280
rect 1632 9220 1636 9276
rect 1636 9220 1692 9276
rect 1692 9220 1696 9276
rect 1632 9216 1696 9220
rect 1712 9276 1776 9280
rect 1712 9220 1716 9276
rect 1716 9220 1772 9276
rect 1772 9220 1776 9276
rect 1712 9216 1776 9220
rect 1792 9276 1856 9280
rect 1792 9220 1796 9276
rect 1796 9220 1852 9276
rect 1852 9220 1856 9276
rect 1792 9216 1856 9220
rect 5552 9276 5616 9280
rect 5552 9220 5556 9276
rect 5556 9220 5612 9276
rect 5612 9220 5616 9276
rect 5552 9216 5616 9220
rect 5632 9276 5696 9280
rect 5632 9220 5636 9276
rect 5636 9220 5692 9276
rect 5692 9220 5696 9276
rect 5632 9216 5696 9220
rect 5712 9276 5776 9280
rect 5712 9220 5716 9276
rect 5716 9220 5772 9276
rect 5772 9220 5776 9276
rect 5712 9216 5776 9220
rect 5792 9276 5856 9280
rect 5792 9220 5796 9276
rect 5796 9220 5852 9276
rect 5852 9220 5856 9276
rect 5792 9216 5856 9220
rect 9552 9276 9616 9280
rect 9552 9220 9556 9276
rect 9556 9220 9612 9276
rect 9612 9220 9616 9276
rect 9552 9216 9616 9220
rect 9632 9276 9696 9280
rect 9632 9220 9636 9276
rect 9636 9220 9692 9276
rect 9692 9220 9696 9276
rect 9632 9216 9696 9220
rect 9712 9276 9776 9280
rect 9712 9220 9716 9276
rect 9716 9220 9772 9276
rect 9772 9220 9776 9276
rect 9712 9216 9776 9220
rect 9792 9276 9856 9280
rect 9792 9220 9796 9276
rect 9796 9220 9852 9276
rect 9852 9220 9856 9276
rect 9792 9216 9856 9220
rect 13552 9276 13616 9280
rect 13552 9220 13556 9276
rect 13556 9220 13612 9276
rect 13612 9220 13616 9276
rect 13552 9216 13616 9220
rect 13632 9276 13696 9280
rect 13632 9220 13636 9276
rect 13636 9220 13692 9276
rect 13692 9220 13696 9276
rect 13632 9216 13696 9220
rect 13712 9276 13776 9280
rect 13712 9220 13716 9276
rect 13716 9220 13772 9276
rect 13772 9220 13776 9276
rect 13712 9216 13776 9220
rect 13792 9276 13856 9280
rect 13792 9220 13796 9276
rect 13796 9220 13852 9276
rect 13852 9220 13856 9276
rect 13792 9216 13856 9220
rect 17552 9276 17616 9280
rect 17552 9220 17556 9276
rect 17556 9220 17612 9276
rect 17612 9220 17616 9276
rect 17552 9216 17616 9220
rect 17632 9276 17696 9280
rect 17632 9220 17636 9276
rect 17636 9220 17692 9276
rect 17692 9220 17696 9276
rect 17632 9216 17696 9220
rect 17712 9276 17776 9280
rect 17712 9220 17716 9276
rect 17716 9220 17772 9276
rect 17772 9220 17776 9276
rect 17712 9216 17776 9220
rect 17792 9276 17856 9280
rect 17792 9220 17796 9276
rect 17796 9220 17852 9276
rect 17852 9220 17856 9276
rect 17792 9216 17856 9220
rect 2212 8732 2276 8736
rect 2212 8676 2216 8732
rect 2216 8676 2272 8732
rect 2272 8676 2276 8732
rect 2212 8672 2276 8676
rect 2292 8732 2356 8736
rect 2292 8676 2296 8732
rect 2296 8676 2352 8732
rect 2352 8676 2356 8732
rect 2292 8672 2356 8676
rect 2372 8732 2436 8736
rect 2372 8676 2376 8732
rect 2376 8676 2432 8732
rect 2432 8676 2436 8732
rect 2372 8672 2436 8676
rect 2452 8732 2516 8736
rect 2452 8676 2456 8732
rect 2456 8676 2512 8732
rect 2512 8676 2516 8732
rect 2452 8672 2516 8676
rect 6212 8732 6276 8736
rect 6212 8676 6216 8732
rect 6216 8676 6272 8732
rect 6272 8676 6276 8732
rect 6212 8672 6276 8676
rect 6292 8732 6356 8736
rect 6292 8676 6296 8732
rect 6296 8676 6352 8732
rect 6352 8676 6356 8732
rect 6292 8672 6356 8676
rect 6372 8732 6436 8736
rect 6372 8676 6376 8732
rect 6376 8676 6432 8732
rect 6432 8676 6436 8732
rect 6372 8672 6436 8676
rect 6452 8732 6516 8736
rect 6452 8676 6456 8732
rect 6456 8676 6512 8732
rect 6512 8676 6516 8732
rect 6452 8672 6516 8676
rect 10212 8732 10276 8736
rect 10212 8676 10216 8732
rect 10216 8676 10272 8732
rect 10272 8676 10276 8732
rect 10212 8672 10276 8676
rect 10292 8732 10356 8736
rect 10292 8676 10296 8732
rect 10296 8676 10352 8732
rect 10352 8676 10356 8732
rect 10292 8672 10356 8676
rect 10372 8732 10436 8736
rect 10372 8676 10376 8732
rect 10376 8676 10432 8732
rect 10432 8676 10436 8732
rect 10372 8672 10436 8676
rect 10452 8732 10516 8736
rect 10452 8676 10456 8732
rect 10456 8676 10512 8732
rect 10512 8676 10516 8732
rect 10452 8672 10516 8676
rect 14212 8732 14276 8736
rect 14212 8676 14216 8732
rect 14216 8676 14272 8732
rect 14272 8676 14276 8732
rect 14212 8672 14276 8676
rect 14292 8732 14356 8736
rect 14292 8676 14296 8732
rect 14296 8676 14352 8732
rect 14352 8676 14356 8732
rect 14292 8672 14356 8676
rect 14372 8732 14436 8736
rect 14372 8676 14376 8732
rect 14376 8676 14432 8732
rect 14432 8676 14436 8732
rect 14372 8672 14436 8676
rect 14452 8732 14516 8736
rect 14452 8676 14456 8732
rect 14456 8676 14512 8732
rect 14512 8676 14516 8732
rect 14452 8672 14516 8676
rect 18212 8732 18276 8736
rect 18212 8676 18216 8732
rect 18216 8676 18272 8732
rect 18272 8676 18276 8732
rect 18212 8672 18276 8676
rect 18292 8732 18356 8736
rect 18292 8676 18296 8732
rect 18296 8676 18352 8732
rect 18352 8676 18356 8732
rect 18292 8672 18356 8676
rect 18372 8732 18436 8736
rect 18372 8676 18376 8732
rect 18376 8676 18432 8732
rect 18432 8676 18436 8732
rect 18372 8672 18436 8676
rect 18452 8732 18516 8736
rect 18452 8676 18456 8732
rect 18456 8676 18512 8732
rect 18512 8676 18516 8732
rect 18452 8672 18516 8676
rect 1552 8188 1616 8192
rect 1552 8132 1556 8188
rect 1556 8132 1612 8188
rect 1612 8132 1616 8188
rect 1552 8128 1616 8132
rect 1632 8188 1696 8192
rect 1632 8132 1636 8188
rect 1636 8132 1692 8188
rect 1692 8132 1696 8188
rect 1632 8128 1696 8132
rect 1712 8188 1776 8192
rect 1712 8132 1716 8188
rect 1716 8132 1772 8188
rect 1772 8132 1776 8188
rect 1712 8128 1776 8132
rect 1792 8188 1856 8192
rect 1792 8132 1796 8188
rect 1796 8132 1852 8188
rect 1852 8132 1856 8188
rect 1792 8128 1856 8132
rect 5552 8188 5616 8192
rect 5552 8132 5556 8188
rect 5556 8132 5612 8188
rect 5612 8132 5616 8188
rect 5552 8128 5616 8132
rect 5632 8188 5696 8192
rect 5632 8132 5636 8188
rect 5636 8132 5692 8188
rect 5692 8132 5696 8188
rect 5632 8128 5696 8132
rect 5712 8188 5776 8192
rect 5712 8132 5716 8188
rect 5716 8132 5772 8188
rect 5772 8132 5776 8188
rect 5712 8128 5776 8132
rect 5792 8188 5856 8192
rect 5792 8132 5796 8188
rect 5796 8132 5852 8188
rect 5852 8132 5856 8188
rect 5792 8128 5856 8132
rect 9552 8188 9616 8192
rect 9552 8132 9556 8188
rect 9556 8132 9612 8188
rect 9612 8132 9616 8188
rect 9552 8128 9616 8132
rect 9632 8188 9696 8192
rect 9632 8132 9636 8188
rect 9636 8132 9692 8188
rect 9692 8132 9696 8188
rect 9632 8128 9696 8132
rect 9712 8188 9776 8192
rect 9712 8132 9716 8188
rect 9716 8132 9772 8188
rect 9772 8132 9776 8188
rect 9712 8128 9776 8132
rect 9792 8188 9856 8192
rect 9792 8132 9796 8188
rect 9796 8132 9852 8188
rect 9852 8132 9856 8188
rect 9792 8128 9856 8132
rect 13552 8188 13616 8192
rect 13552 8132 13556 8188
rect 13556 8132 13612 8188
rect 13612 8132 13616 8188
rect 13552 8128 13616 8132
rect 13632 8188 13696 8192
rect 13632 8132 13636 8188
rect 13636 8132 13692 8188
rect 13692 8132 13696 8188
rect 13632 8128 13696 8132
rect 13712 8188 13776 8192
rect 13712 8132 13716 8188
rect 13716 8132 13772 8188
rect 13772 8132 13776 8188
rect 13712 8128 13776 8132
rect 13792 8188 13856 8192
rect 13792 8132 13796 8188
rect 13796 8132 13852 8188
rect 13852 8132 13856 8188
rect 13792 8128 13856 8132
rect 17552 8188 17616 8192
rect 17552 8132 17556 8188
rect 17556 8132 17612 8188
rect 17612 8132 17616 8188
rect 17552 8128 17616 8132
rect 17632 8188 17696 8192
rect 17632 8132 17636 8188
rect 17636 8132 17692 8188
rect 17692 8132 17696 8188
rect 17632 8128 17696 8132
rect 17712 8188 17776 8192
rect 17712 8132 17716 8188
rect 17716 8132 17772 8188
rect 17772 8132 17776 8188
rect 17712 8128 17776 8132
rect 17792 8188 17856 8192
rect 17792 8132 17796 8188
rect 17796 8132 17852 8188
rect 17852 8132 17856 8188
rect 17792 8128 17856 8132
rect 2212 7644 2276 7648
rect 2212 7588 2216 7644
rect 2216 7588 2272 7644
rect 2272 7588 2276 7644
rect 2212 7584 2276 7588
rect 2292 7644 2356 7648
rect 2292 7588 2296 7644
rect 2296 7588 2352 7644
rect 2352 7588 2356 7644
rect 2292 7584 2356 7588
rect 2372 7644 2436 7648
rect 2372 7588 2376 7644
rect 2376 7588 2432 7644
rect 2432 7588 2436 7644
rect 2372 7584 2436 7588
rect 2452 7644 2516 7648
rect 2452 7588 2456 7644
rect 2456 7588 2512 7644
rect 2512 7588 2516 7644
rect 2452 7584 2516 7588
rect 6212 7644 6276 7648
rect 6212 7588 6216 7644
rect 6216 7588 6272 7644
rect 6272 7588 6276 7644
rect 6212 7584 6276 7588
rect 6292 7644 6356 7648
rect 6292 7588 6296 7644
rect 6296 7588 6352 7644
rect 6352 7588 6356 7644
rect 6292 7584 6356 7588
rect 6372 7644 6436 7648
rect 6372 7588 6376 7644
rect 6376 7588 6432 7644
rect 6432 7588 6436 7644
rect 6372 7584 6436 7588
rect 6452 7644 6516 7648
rect 6452 7588 6456 7644
rect 6456 7588 6512 7644
rect 6512 7588 6516 7644
rect 6452 7584 6516 7588
rect 10212 7644 10276 7648
rect 10212 7588 10216 7644
rect 10216 7588 10272 7644
rect 10272 7588 10276 7644
rect 10212 7584 10276 7588
rect 10292 7644 10356 7648
rect 10292 7588 10296 7644
rect 10296 7588 10352 7644
rect 10352 7588 10356 7644
rect 10292 7584 10356 7588
rect 10372 7644 10436 7648
rect 10372 7588 10376 7644
rect 10376 7588 10432 7644
rect 10432 7588 10436 7644
rect 10372 7584 10436 7588
rect 10452 7644 10516 7648
rect 10452 7588 10456 7644
rect 10456 7588 10512 7644
rect 10512 7588 10516 7644
rect 10452 7584 10516 7588
rect 14212 7644 14276 7648
rect 14212 7588 14216 7644
rect 14216 7588 14272 7644
rect 14272 7588 14276 7644
rect 14212 7584 14276 7588
rect 14292 7644 14356 7648
rect 14292 7588 14296 7644
rect 14296 7588 14352 7644
rect 14352 7588 14356 7644
rect 14292 7584 14356 7588
rect 14372 7644 14436 7648
rect 14372 7588 14376 7644
rect 14376 7588 14432 7644
rect 14432 7588 14436 7644
rect 14372 7584 14436 7588
rect 14452 7644 14516 7648
rect 14452 7588 14456 7644
rect 14456 7588 14512 7644
rect 14512 7588 14516 7644
rect 14452 7584 14516 7588
rect 18212 7644 18276 7648
rect 18212 7588 18216 7644
rect 18216 7588 18272 7644
rect 18272 7588 18276 7644
rect 18212 7584 18276 7588
rect 18292 7644 18356 7648
rect 18292 7588 18296 7644
rect 18296 7588 18352 7644
rect 18352 7588 18356 7644
rect 18292 7584 18356 7588
rect 18372 7644 18436 7648
rect 18372 7588 18376 7644
rect 18376 7588 18432 7644
rect 18432 7588 18436 7644
rect 18372 7584 18436 7588
rect 18452 7644 18516 7648
rect 18452 7588 18456 7644
rect 18456 7588 18512 7644
rect 18512 7588 18516 7644
rect 18452 7584 18516 7588
rect 1552 7100 1616 7104
rect 1552 7044 1556 7100
rect 1556 7044 1612 7100
rect 1612 7044 1616 7100
rect 1552 7040 1616 7044
rect 1632 7100 1696 7104
rect 1632 7044 1636 7100
rect 1636 7044 1692 7100
rect 1692 7044 1696 7100
rect 1632 7040 1696 7044
rect 1712 7100 1776 7104
rect 1712 7044 1716 7100
rect 1716 7044 1772 7100
rect 1772 7044 1776 7100
rect 1712 7040 1776 7044
rect 1792 7100 1856 7104
rect 1792 7044 1796 7100
rect 1796 7044 1852 7100
rect 1852 7044 1856 7100
rect 1792 7040 1856 7044
rect 5552 7100 5616 7104
rect 5552 7044 5556 7100
rect 5556 7044 5612 7100
rect 5612 7044 5616 7100
rect 5552 7040 5616 7044
rect 5632 7100 5696 7104
rect 5632 7044 5636 7100
rect 5636 7044 5692 7100
rect 5692 7044 5696 7100
rect 5632 7040 5696 7044
rect 5712 7100 5776 7104
rect 5712 7044 5716 7100
rect 5716 7044 5772 7100
rect 5772 7044 5776 7100
rect 5712 7040 5776 7044
rect 5792 7100 5856 7104
rect 5792 7044 5796 7100
rect 5796 7044 5852 7100
rect 5852 7044 5856 7100
rect 5792 7040 5856 7044
rect 9552 7100 9616 7104
rect 9552 7044 9556 7100
rect 9556 7044 9612 7100
rect 9612 7044 9616 7100
rect 9552 7040 9616 7044
rect 9632 7100 9696 7104
rect 9632 7044 9636 7100
rect 9636 7044 9692 7100
rect 9692 7044 9696 7100
rect 9632 7040 9696 7044
rect 9712 7100 9776 7104
rect 9712 7044 9716 7100
rect 9716 7044 9772 7100
rect 9772 7044 9776 7100
rect 9712 7040 9776 7044
rect 9792 7100 9856 7104
rect 9792 7044 9796 7100
rect 9796 7044 9852 7100
rect 9852 7044 9856 7100
rect 9792 7040 9856 7044
rect 13552 7100 13616 7104
rect 13552 7044 13556 7100
rect 13556 7044 13612 7100
rect 13612 7044 13616 7100
rect 13552 7040 13616 7044
rect 13632 7100 13696 7104
rect 13632 7044 13636 7100
rect 13636 7044 13692 7100
rect 13692 7044 13696 7100
rect 13632 7040 13696 7044
rect 13712 7100 13776 7104
rect 13712 7044 13716 7100
rect 13716 7044 13772 7100
rect 13772 7044 13776 7100
rect 13712 7040 13776 7044
rect 13792 7100 13856 7104
rect 13792 7044 13796 7100
rect 13796 7044 13852 7100
rect 13852 7044 13856 7100
rect 13792 7040 13856 7044
rect 17552 7100 17616 7104
rect 17552 7044 17556 7100
rect 17556 7044 17612 7100
rect 17612 7044 17616 7100
rect 17552 7040 17616 7044
rect 17632 7100 17696 7104
rect 17632 7044 17636 7100
rect 17636 7044 17692 7100
rect 17692 7044 17696 7100
rect 17632 7040 17696 7044
rect 17712 7100 17776 7104
rect 17712 7044 17716 7100
rect 17716 7044 17772 7100
rect 17772 7044 17776 7100
rect 17712 7040 17776 7044
rect 17792 7100 17856 7104
rect 17792 7044 17796 7100
rect 17796 7044 17852 7100
rect 17852 7044 17856 7100
rect 17792 7040 17856 7044
rect 2212 6556 2276 6560
rect 2212 6500 2216 6556
rect 2216 6500 2272 6556
rect 2272 6500 2276 6556
rect 2212 6496 2276 6500
rect 2292 6556 2356 6560
rect 2292 6500 2296 6556
rect 2296 6500 2352 6556
rect 2352 6500 2356 6556
rect 2292 6496 2356 6500
rect 2372 6556 2436 6560
rect 2372 6500 2376 6556
rect 2376 6500 2432 6556
rect 2432 6500 2436 6556
rect 2372 6496 2436 6500
rect 2452 6556 2516 6560
rect 2452 6500 2456 6556
rect 2456 6500 2512 6556
rect 2512 6500 2516 6556
rect 2452 6496 2516 6500
rect 6212 6556 6276 6560
rect 6212 6500 6216 6556
rect 6216 6500 6272 6556
rect 6272 6500 6276 6556
rect 6212 6496 6276 6500
rect 6292 6556 6356 6560
rect 6292 6500 6296 6556
rect 6296 6500 6352 6556
rect 6352 6500 6356 6556
rect 6292 6496 6356 6500
rect 6372 6556 6436 6560
rect 6372 6500 6376 6556
rect 6376 6500 6432 6556
rect 6432 6500 6436 6556
rect 6372 6496 6436 6500
rect 6452 6556 6516 6560
rect 6452 6500 6456 6556
rect 6456 6500 6512 6556
rect 6512 6500 6516 6556
rect 6452 6496 6516 6500
rect 10212 6556 10276 6560
rect 10212 6500 10216 6556
rect 10216 6500 10272 6556
rect 10272 6500 10276 6556
rect 10212 6496 10276 6500
rect 10292 6556 10356 6560
rect 10292 6500 10296 6556
rect 10296 6500 10352 6556
rect 10352 6500 10356 6556
rect 10292 6496 10356 6500
rect 10372 6556 10436 6560
rect 10372 6500 10376 6556
rect 10376 6500 10432 6556
rect 10432 6500 10436 6556
rect 10372 6496 10436 6500
rect 10452 6556 10516 6560
rect 10452 6500 10456 6556
rect 10456 6500 10512 6556
rect 10512 6500 10516 6556
rect 10452 6496 10516 6500
rect 14212 6556 14276 6560
rect 14212 6500 14216 6556
rect 14216 6500 14272 6556
rect 14272 6500 14276 6556
rect 14212 6496 14276 6500
rect 14292 6556 14356 6560
rect 14292 6500 14296 6556
rect 14296 6500 14352 6556
rect 14352 6500 14356 6556
rect 14292 6496 14356 6500
rect 14372 6556 14436 6560
rect 14372 6500 14376 6556
rect 14376 6500 14432 6556
rect 14432 6500 14436 6556
rect 14372 6496 14436 6500
rect 14452 6556 14516 6560
rect 14452 6500 14456 6556
rect 14456 6500 14512 6556
rect 14512 6500 14516 6556
rect 14452 6496 14516 6500
rect 18212 6556 18276 6560
rect 18212 6500 18216 6556
rect 18216 6500 18272 6556
rect 18272 6500 18276 6556
rect 18212 6496 18276 6500
rect 18292 6556 18356 6560
rect 18292 6500 18296 6556
rect 18296 6500 18352 6556
rect 18352 6500 18356 6556
rect 18292 6496 18356 6500
rect 18372 6556 18436 6560
rect 18372 6500 18376 6556
rect 18376 6500 18432 6556
rect 18432 6500 18436 6556
rect 18372 6496 18436 6500
rect 18452 6556 18516 6560
rect 18452 6500 18456 6556
rect 18456 6500 18512 6556
rect 18512 6500 18516 6556
rect 18452 6496 18516 6500
rect 1552 6012 1616 6016
rect 1552 5956 1556 6012
rect 1556 5956 1612 6012
rect 1612 5956 1616 6012
rect 1552 5952 1616 5956
rect 1632 6012 1696 6016
rect 1632 5956 1636 6012
rect 1636 5956 1692 6012
rect 1692 5956 1696 6012
rect 1632 5952 1696 5956
rect 1712 6012 1776 6016
rect 1712 5956 1716 6012
rect 1716 5956 1772 6012
rect 1772 5956 1776 6012
rect 1712 5952 1776 5956
rect 1792 6012 1856 6016
rect 1792 5956 1796 6012
rect 1796 5956 1852 6012
rect 1852 5956 1856 6012
rect 1792 5952 1856 5956
rect 5552 6012 5616 6016
rect 5552 5956 5556 6012
rect 5556 5956 5612 6012
rect 5612 5956 5616 6012
rect 5552 5952 5616 5956
rect 5632 6012 5696 6016
rect 5632 5956 5636 6012
rect 5636 5956 5692 6012
rect 5692 5956 5696 6012
rect 5632 5952 5696 5956
rect 5712 6012 5776 6016
rect 5712 5956 5716 6012
rect 5716 5956 5772 6012
rect 5772 5956 5776 6012
rect 5712 5952 5776 5956
rect 5792 6012 5856 6016
rect 5792 5956 5796 6012
rect 5796 5956 5852 6012
rect 5852 5956 5856 6012
rect 5792 5952 5856 5956
rect 9552 6012 9616 6016
rect 9552 5956 9556 6012
rect 9556 5956 9612 6012
rect 9612 5956 9616 6012
rect 9552 5952 9616 5956
rect 9632 6012 9696 6016
rect 9632 5956 9636 6012
rect 9636 5956 9692 6012
rect 9692 5956 9696 6012
rect 9632 5952 9696 5956
rect 9712 6012 9776 6016
rect 9712 5956 9716 6012
rect 9716 5956 9772 6012
rect 9772 5956 9776 6012
rect 9712 5952 9776 5956
rect 9792 6012 9856 6016
rect 9792 5956 9796 6012
rect 9796 5956 9852 6012
rect 9852 5956 9856 6012
rect 9792 5952 9856 5956
rect 13552 6012 13616 6016
rect 13552 5956 13556 6012
rect 13556 5956 13612 6012
rect 13612 5956 13616 6012
rect 13552 5952 13616 5956
rect 13632 6012 13696 6016
rect 13632 5956 13636 6012
rect 13636 5956 13692 6012
rect 13692 5956 13696 6012
rect 13632 5952 13696 5956
rect 13712 6012 13776 6016
rect 13712 5956 13716 6012
rect 13716 5956 13772 6012
rect 13772 5956 13776 6012
rect 13712 5952 13776 5956
rect 13792 6012 13856 6016
rect 13792 5956 13796 6012
rect 13796 5956 13852 6012
rect 13852 5956 13856 6012
rect 13792 5952 13856 5956
rect 17552 6012 17616 6016
rect 17552 5956 17556 6012
rect 17556 5956 17612 6012
rect 17612 5956 17616 6012
rect 17552 5952 17616 5956
rect 17632 6012 17696 6016
rect 17632 5956 17636 6012
rect 17636 5956 17692 6012
rect 17692 5956 17696 6012
rect 17632 5952 17696 5956
rect 17712 6012 17776 6016
rect 17712 5956 17716 6012
rect 17716 5956 17772 6012
rect 17772 5956 17776 6012
rect 17712 5952 17776 5956
rect 17792 6012 17856 6016
rect 17792 5956 17796 6012
rect 17796 5956 17852 6012
rect 17852 5956 17856 6012
rect 17792 5952 17856 5956
rect 2212 5468 2276 5472
rect 2212 5412 2216 5468
rect 2216 5412 2272 5468
rect 2272 5412 2276 5468
rect 2212 5408 2276 5412
rect 2292 5468 2356 5472
rect 2292 5412 2296 5468
rect 2296 5412 2352 5468
rect 2352 5412 2356 5468
rect 2292 5408 2356 5412
rect 2372 5468 2436 5472
rect 2372 5412 2376 5468
rect 2376 5412 2432 5468
rect 2432 5412 2436 5468
rect 2372 5408 2436 5412
rect 2452 5468 2516 5472
rect 2452 5412 2456 5468
rect 2456 5412 2512 5468
rect 2512 5412 2516 5468
rect 2452 5408 2516 5412
rect 6212 5468 6276 5472
rect 6212 5412 6216 5468
rect 6216 5412 6272 5468
rect 6272 5412 6276 5468
rect 6212 5408 6276 5412
rect 6292 5468 6356 5472
rect 6292 5412 6296 5468
rect 6296 5412 6352 5468
rect 6352 5412 6356 5468
rect 6292 5408 6356 5412
rect 6372 5468 6436 5472
rect 6372 5412 6376 5468
rect 6376 5412 6432 5468
rect 6432 5412 6436 5468
rect 6372 5408 6436 5412
rect 6452 5468 6516 5472
rect 6452 5412 6456 5468
rect 6456 5412 6512 5468
rect 6512 5412 6516 5468
rect 6452 5408 6516 5412
rect 10212 5468 10276 5472
rect 10212 5412 10216 5468
rect 10216 5412 10272 5468
rect 10272 5412 10276 5468
rect 10212 5408 10276 5412
rect 10292 5468 10356 5472
rect 10292 5412 10296 5468
rect 10296 5412 10352 5468
rect 10352 5412 10356 5468
rect 10292 5408 10356 5412
rect 10372 5468 10436 5472
rect 10372 5412 10376 5468
rect 10376 5412 10432 5468
rect 10432 5412 10436 5468
rect 10372 5408 10436 5412
rect 10452 5468 10516 5472
rect 10452 5412 10456 5468
rect 10456 5412 10512 5468
rect 10512 5412 10516 5468
rect 10452 5408 10516 5412
rect 14212 5468 14276 5472
rect 14212 5412 14216 5468
rect 14216 5412 14272 5468
rect 14272 5412 14276 5468
rect 14212 5408 14276 5412
rect 14292 5468 14356 5472
rect 14292 5412 14296 5468
rect 14296 5412 14352 5468
rect 14352 5412 14356 5468
rect 14292 5408 14356 5412
rect 14372 5468 14436 5472
rect 14372 5412 14376 5468
rect 14376 5412 14432 5468
rect 14432 5412 14436 5468
rect 14372 5408 14436 5412
rect 14452 5468 14516 5472
rect 14452 5412 14456 5468
rect 14456 5412 14512 5468
rect 14512 5412 14516 5468
rect 14452 5408 14516 5412
rect 18212 5468 18276 5472
rect 18212 5412 18216 5468
rect 18216 5412 18272 5468
rect 18272 5412 18276 5468
rect 18212 5408 18276 5412
rect 18292 5468 18356 5472
rect 18292 5412 18296 5468
rect 18296 5412 18352 5468
rect 18352 5412 18356 5468
rect 18292 5408 18356 5412
rect 18372 5468 18436 5472
rect 18372 5412 18376 5468
rect 18376 5412 18432 5468
rect 18432 5412 18436 5468
rect 18372 5408 18436 5412
rect 18452 5468 18516 5472
rect 18452 5412 18456 5468
rect 18456 5412 18512 5468
rect 18512 5412 18516 5468
rect 18452 5408 18516 5412
rect 1552 4924 1616 4928
rect 1552 4868 1556 4924
rect 1556 4868 1612 4924
rect 1612 4868 1616 4924
rect 1552 4864 1616 4868
rect 1632 4924 1696 4928
rect 1632 4868 1636 4924
rect 1636 4868 1692 4924
rect 1692 4868 1696 4924
rect 1632 4864 1696 4868
rect 1712 4924 1776 4928
rect 1712 4868 1716 4924
rect 1716 4868 1772 4924
rect 1772 4868 1776 4924
rect 1712 4864 1776 4868
rect 1792 4924 1856 4928
rect 1792 4868 1796 4924
rect 1796 4868 1852 4924
rect 1852 4868 1856 4924
rect 1792 4864 1856 4868
rect 5552 4924 5616 4928
rect 5552 4868 5556 4924
rect 5556 4868 5612 4924
rect 5612 4868 5616 4924
rect 5552 4864 5616 4868
rect 5632 4924 5696 4928
rect 5632 4868 5636 4924
rect 5636 4868 5692 4924
rect 5692 4868 5696 4924
rect 5632 4864 5696 4868
rect 5712 4924 5776 4928
rect 5712 4868 5716 4924
rect 5716 4868 5772 4924
rect 5772 4868 5776 4924
rect 5712 4864 5776 4868
rect 5792 4924 5856 4928
rect 5792 4868 5796 4924
rect 5796 4868 5852 4924
rect 5852 4868 5856 4924
rect 5792 4864 5856 4868
rect 9552 4924 9616 4928
rect 9552 4868 9556 4924
rect 9556 4868 9612 4924
rect 9612 4868 9616 4924
rect 9552 4864 9616 4868
rect 9632 4924 9696 4928
rect 9632 4868 9636 4924
rect 9636 4868 9692 4924
rect 9692 4868 9696 4924
rect 9632 4864 9696 4868
rect 9712 4924 9776 4928
rect 9712 4868 9716 4924
rect 9716 4868 9772 4924
rect 9772 4868 9776 4924
rect 9712 4864 9776 4868
rect 9792 4924 9856 4928
rect 9792 4868 9796 4924
rect 9796 4868 9852 4924
rect 9852 4868 9856 4924
rect 9792 4864 9856 4868
rect 13552 4924 13616 4928
rect 13552 4868 13556 4924
rect 13556 4868 13612 4924
rect 13612 4868 13616 4924
rect 13552 4864 13616 4868
rect 13632 4924 13696 4928
rect 13632 4868 13636 4924
rect 13636 4868 13692 4924
rect 13692 4868 13696 4924
rect 13632 4864 13696 4868
rect 13712 4924 13776 4928
rect 13712 4868 13716 4924
rect 13716 4868 13772 4924
rect 13772 4868 13776 4924
rect 13712 4864 13776 4868
rect 13792 4924 13856 4928
rect 13792 4868 13796 4924
rect 13796 4868 13852 4924
rect 13852 4868 13856 4924
rect 13792 4864 13856 4868
rect 17552 4924 17616 4928
rect 17552 4868 17556 4924
rect 17556 4868 17612 4924
rect 17612 4868 17616 4924
rect 17552 4864 17616 4868
rect 17632 4924 17696 4928
rect 17632 4868 17636 4924
rect 17636 4868 17692 4924
rect 17692 4868 17696 4924
rect 17632 4864 17696 4868
rect 17712 4924 17776 4928
rect 17712 4868 17716 4924
rect 17716 4868 17772 4924
rect 17772 4868 17776 4924
rect 17712 4864 17776 4868
rect 17792 4924 17856 4928
rect 17792 4868 17796 4924
rect 17796 4868 17852 4924
rect 17852 4868 17856 4924
rect 17792 4864 17856 4868
rect 2212 4380 2276 4384
rect 2212 4324 2216 4380
rect 2216 4324 2272 4380
rect 2272 4324 2276 4380
rect 2212 4320 2276 4324
rect 2292 4380 2356 4384
rect 2292 4324 2296 4380
rect 2296 4324 2352 4380
rect 2352 4324 2356 4380
rect 2292 4320 2356 4324
rect 2372 4380 2436 4384
rect 2372 4324 2376 4380
rect 2376 4324 2432 4380
rect 2432 4324 2436 4380
rect 2372 4320 2436 4324
rect 2452 4380 2516 4384
rect 2452 4324 2456 4380
rect 2456 4324 2512 4380
rect 2512 4324 2516 4380
rect 2452 4320 2516 4324
rect 6212 4380 6276 4384
rect 6212 4324 6216 4380
rect 6216 4324 6272 4380
rect 6272 4324 6276 4380
rect 6212 4320 6276 4324
rect 6292 4380 6356 4384
rect 6292 4324 6296 4380
rect 6296 4324 6352 4380
rect 6352 4324 6356 4380
rect 6292 4320 6356 4324
rect 6372 4380 6436 4384
rect 6372 4324 6376 4380
rect 6376 4324 6432 4380
rect 6432 4324 6436 4380
rect 6372 4320 6436 4324
rect 6452 4380 6516 4384
rect 6452 4324 6456 4380
rect 6456 4324 6512 4380
rect 6512 4324 6516 4380
rect 6452 4320 6516 4324
rect 10212 4380 10276 4384
rect 10212 4324 10216 4380
rect 10216 4324 10272 4380
rect 10272 4324 10276 4380
rect 10212 4320 10276 4324
rect 10292 4380 10356 4384
rect 10292 4324 10296 4380
rect 10296 4324 10352 4380
rect 10352 4324 10356 4380
rect 10292 4320 10356 4324
rect 10372 4380 10436 4384
rect 10372 4324 10376 4380
rect 10376 4324 10432 4380
rect 10432 4324 10436 4380
rect 10372 4320 10436 4324
rect 10452 4380 10516 4384
rect 10452 4324 10456 4380
rect 10456 4324 10512 4380
rect 10512 4324 10516 4380
rect 10452 4320 10516 4324
rect 14212 4380 14276 4384
rect 14212 4324 14216 4380
rect 14216 4324 14272 4380
rect 14272 4324 14276 4380
rect 14212 4320 14276 4324
rect 14292 4380 14356 4384
rect 14292 4324 14296 4380
rect 14296 4324 14352 4380
rect 14352 4324 14356 4380
rect 14292 4320 14356 4324
rect 14372 4380 14436 4384
rect 14372 4324 14376 4380
rect 14376 4324 14432 4380
rect 14432 4324 14436 4380
rect 14372 4320 14436 4324
rect 14452 4380 14516 4384
rect 14452 4324 14456 4380
rect 14456 4324 14512 4380
rect 14512 4324 14516 4380
rect 14452 4320 14516 4324
rect 18212 4380 18276 4384
rect 18212 4324 18216 4380
rect 18216 4324 18272 4380
rect 18272 4324 18276 4380
rect 18212 4320 18276 4324
rect 18292 4380 18356 4384
rect 18292 4324 18296 4380
rect 18296 4324 18352 4380
rect 18352 4324 18356 4380
rect 18292 4320 18356 4324
rect 18372 4380 18436 4384
rect 18372 4324 18376 4380
rect 18376 4324 18432 4380
rect 18432 4324 18436 4380
rect 18372 4320 18436 4324
rect 18452 4380 18516 4384
rect 18452 4324 18456 4380
rect 18456 4324 18512 4380
rect 18512 4324 18516 4380
rect 18452 4320 18516 4324
rect 1552 3836 1616 3840
rect 1552 3780 1556 3836
rect 1556 3780 1612 3836
rect 1612 3780 1616 3836
rect 1552 3776 1616 3780
rect 1632 3836 1696 3840
rect 1632 3780 1636 3836
rect 1636 3780 1692 3836
rect 1692 3780 1696 3836
rect 1632 3776 1696 3780
rect 1712 3836 1776 3840
rect 1712 3780 1716 3836
rect 1716 3780 1772 3836
rect 1772 3780 1776 3836
rect 1712 3776 1776 3780
rect 1792 3836 1856 3840
rect 1792 3780 1796 3836
rect 1796 3780 1852 3836
rect 1852 3780 1856 3836
rect 1792 3776 1856 3780
rect 5552 3836 5616 3840
rect 5552 3780 5556 3836
rect 5556 3780 5612 3836
rect 5612 3780 5616 3836
rect 5552 3776 5616 3780
rect 5632 3836 5696 3840
rect 5632 3780 5636 3836
rect 5636 3780 5692 3836
rect 5692 3780 5696 3836
rect 5632 3776 5696 3780
rect 5712 3836 5776 3840
rect 5712 3780 5716 3836
rect 5716 3780 5772 3836
rect 5772 3780 5776 3836
rect 5712 3776 5776 3780
rect 5792 3836 5856 3840
rect 5792 3780 5796 3836
rect 5796 3780 5852 3836
rect 5852 3780 5856 3836
rect 5792 3776 5856 3780
rect 9552 3836 9616 3840
rect 9552 3780 9556 3836
rect 9556 3780 9612 3836
rect 9612 3780 9616 3836
rect 9552 3776 9616 3780
rect 9632 3836 9696 3840
rect 9632 3780 9636 3836
rect 9636 3780 9692 3836
rect 9692 3780 9696 3836
rect 9632 3776 9696 3780
rect 9712 3836 9776 3840
rect 9712 3780 9716 3836
rect 9716 3780 9772 3836
rect 9772 3780 9776 3836
rect 9712 3776 9776 3780
rect 9792 3836 9856 3840
rect 9792 3780 9796 3836
rect 9796 3780 9852 3836
rect 9852 3780 9856 3836
rect 9792 3776 9856 3780
rect 13552 3836 13616 3840
rect 13552 3780 13556 3836
rect 13556 3780 13612 3836
rect 13612 3780 13616 3836
rect 13552 3776 13616 3780
rect 13632 3836 13696 3840
rect 13632 3780 13636 3836
rect 13636 3780 13692 3836
rect 13692 3780 13696 3836
rect 13632 3776 13696 3780
rect 13712 3836 13776 3840
rect 13712 3780 13716 3836
rect 13716 3780 13772 3836
rect 13772 3780 13776 3836
rect 13712 3776 13776 3780
rect 13792 3836 13856 3840
rect 13792 3780 13796 3836
rect 13796 3780 13852 3836
rect 13852 3780 13856 3836
rect 13792 3776 13856 3780
rect 17552 3836 17616 3840
rect 17552 3780 17556 3836
rect 17556 3780 17612 3836
rect 17612 3780 17616 3836
rect 17552 3776 17616 3780
rect 17632 3836 17696 3840
rect 17632 3780 17636 3836
rect 17636 3780 17692 3836
rect 17692 3780 17696 3836
rect 17632 3776 17696 3780
rect 17712 3836 17776 3840
rect 17712 3780 17716 3836
rect 17716 3780 17772 3836
rect 17772 3780 17776 3836
rect 17712 3776 17776 3780
rect 17792 3836 17856 3840
rect 17792 3780 17796 3836
rect 17796 3780 17852 3836
rect 17852 3780 17856 3836
rect 17792 3776 17856 3780
rect 2212 3292 2276 3296
rect 2212 3236 2216 3292
rect 2216 3236 2272 3292
rect 2272 3236 2276 3292
rect 2212 3232 2276 3236
rect 2292 3292 2356 3296
rect 2292 3236 2296 3292
rect 2296 3236 2352 3292
rect 2352 3236 2356 3292
rect 2292 3232 2356 3236
rect 2372 3292 2436 3296
rect 2372 3236 2376 3292
rect 2376 3236 2432 3292
rect 2432 3236 2436 3292
rect 2372 3232 2436 3236
rect 2452 3292 2516 3296
rect 2452 3236 2456 3292
rect 2456 3236 2512 3292
rect 2512 3236 2516 3292
rect 2452 3232 2516 3236
rect 6212 3292 6276 3296
rect 6212 3236 6216 3292
rect 6216 3236 6272 3292
rect 6272 3236 6276 3292
rect 6212 3232 6276 3236
rect 6292 3292 6356 3296
rect 6292 3236 6296 3292
rect 6296 3236 6352 3292
rect 6352 3236 6356 3292
rect 6292 3232 6356 3236
rect 6372 3292 6436 3296
rect 6372 3236 6376 3292
rect 6376 3236 6432 3292
rect 6432 3236 6436 3292
rect 6372 3232 6436 3236
rect 6452 3292 6516 3296
rect 6452 3236 6456 3292
rect 6456 3236 6512 3292
rect 6512 3236 6516 3292
rect 6452 3232 6516 3236
rect 10212 3292 10276 3296
rect 10212 3236 10216 3292
rect 10216 3236 10272 3292
rect 10272 3236 10276 3292
rect 10212 3232 10276 3236
rect 10292 3292 10356 3296
rect 10292 3236 10296 3292
rect 10296 3236 10352 3292
rect 10352 3236 10356 3292
rect 10292 3232 10356 3236
rect 10372 3292 10436 3296
rect 10372 3236 10376 3292
rect 10376 3236 10432 3292
rect 10432 3236 10436 3292
rect 10372 3232 10436 3236
rect 10452 3292 10516 3296
rect 10452 3236 10456 3292
rect 10456 3236 10512 3292
rect 10512 3236 10516 3292
rect 10452 3232 10516 3236
rect 14212 3292 14276 3296
rect 14212 3236 14216 3292
rect 14216 3236 14272 3292
rect 14272 3236 14276 3292
rect 14212 3232 14276 3236
rect 14292 3292 14356 3296
rect 14292 3236 14296 3292
rect 14296 3236 14352 3292
rect 14352 3236 14356 3292
rect 14292 3232 14356 3236
rect 14372 3292 14436 3296
rect 14372 3236 14376 3292
rect 14376 3236 14432 3292
rect 14432 3236 14436 3292
rect 14372 3232 14436 3236
rect 14452 3292 14516 3296
rect 14452 3236 14456 3292
rect 14456 3236 14512 3292
rect 14512 3236 14516 3292
rect 14452 3232 14516 3236
rect 18212 3292 18276 3296
rect 18212 3236 18216 3292
rect 18216 3236 18272 3292
rect 18272 3236 18276 3292
rect 18212 3232 18276 3236
rect 18292 3292 18356 3296
rect 18292 3236 18296 3292
rect 18296 3236 18352 3292
rect 18352 3236 18356 3292
rect 18292 3232 18356 3236
rect 18372 3292 18436 3296
rect 18372 3236 18376 3292
rect 18376 3236 18432 3292
rect 18432 3236 18436 3292
rect 18372 3232 18436 3236
rect 18452 3292 18516 3296
rect 18452 3236 18456 3292
rect 18456 3236 18512 3292
rect 18512 3236 18516 3292
rect 18452 3232 18516 3236
rect 1552 2748 1616 2752
rect 1552 2692 1556 2748
rect 1556 2692 1612 2748
rect 1612 2692 1616 2748
rect 1552 2688 1616 2692
rect 1632 2748 1696 2752
rect 1632 2692 1636 2748
rect 1636 2692 1692 2748
rect 1692 2692 1696 2748
rect 1632 2688 1696 2692
rect 1712 2748 1776 2752
rect 1712 2692 1716 2748
rect 1716 2692 1772 2748
rect 1772 2692 1776 2748
rect 1712 2688 1776 2692
rect 1792 2748 1856 2752
rect 1792 2692 1796 2748
rect 1796 2692 1852 2748
rect 1852 2692 1856 2748
rect 1792 2688 1856 2692
rect 5552 2748 5616 2752
rect 5552 2692 5556 2748
rect 5556 2692 5612 2748
rect 5612 2692 5616 2748
rect 5552 2688 5616 2692
rect 5632 2748 5696 2752
rect 5632 2692 5636 2748
rect 5636 2692 5692 2748
rect 5692 2692 5696 2748
rect 5632 2688 5696 2692
rect 5712 2748 5776 2752
rect 5712 2692 5716 2748
rect 5716 2692 5772 2748
rect 5772 2692 5776 2748
rect 5712 2688 5776 2692
rect 5792 2748 5856 2752
rect 5792 2692 5796 2748
rect 5796 2692 5852 2748
rect 5852 2692 5856 2748
rect 5792 2688 5856 2692
rect 9552 2748 9616 2752
rect 9552 2692 9556 2748
rect 9556 2692 9612 2748
rect 9612 2692 9616 2748
rect 9552 2688 9616 2692
rect 9632 2748 9696 2752
rect 9632 2692 9636 2748
rect 9636 2692 9692 2748
rect 9692 2692 9696 2748
rect 9632 2688 9696 2692
rect 9712 2748 9776 2752
rect 9712 2692 9716 2748
rect 9716 2692 9772 2748
rect 9772 2692 9776 2748
rect 9712 2688 9776 2692
rect 9792 2748 9856 2752
rect 9792 2692 9796 2748
rect 9796 2692 9852 2748
rect 9852 2692 9856 2748
rect 9792 2688 9856 2692
rect 13552 2748 13616 2752
rect 13552 2692 13556 2748
rect 13556 2692 13612 2748
rect 13612 2692 13616 2748
rect 13552 2688 13616 2692
rect 13632 2748 13696 2752
rect 13632 2692 13636 2748
rect 13636 2692 13692 2748
rect 13692 2692 13696 2748
rect 13632 2688 13696 2692
rect 13712 2748 13776 2752
rect 13712 2692 13716 2748
rect 13716 2692 13772 2748
rect 13772 2692 13776 2748
rect 13712 2688 13776 2692
rect 13792 2748 13856 2752
rect 13792 2692 13796 2748
rect 13796 2692 13852 2748
rect 13852 2692 13856 2748
rect 13792 2688 13856 2692
rect 17552 2748 17616 2752
rect 17552 2692 17556 2748
rect 17556 2692 17612 2748
rect 17612 2692 17616 2748
rect 17552 2688 17616 2692
rect 17632 2748 17696 2752
rect 17632 2692 17636 2748
rect 17636 2692 17692 2748
rect 17692 2692 17696 2748
rect 17632 2688 17696 2692
rect 17712 2748 17776 2752
rect 17712 2692 17716 2748
rect 17716 2692 17772 2748
rect 17772 2692 17776 2748
rect 17712 2688 17776 2692
rect 17792 2748 17856 2752
rect 17792 2692 17796 2748
rect 17796 2692 17852 2748
rect 17852 2692 17856 2748
rect 17792 2688 17856 2692
rect 2212 2204 2276 2208
rect 2212 2148 2216 2204
rect 2216 2148 2272 2204
rect 2272 2148 2276 2204
rect 2212 2144 2276 2148
rect 2292 2204 2356 2208
rect 2292 2148 2296 2204
rect 2296 2148 2352 2204
rect 2352 2148 2356 2204
rect 2292 2144 2356 2148
rect 2372 2204 2436 2208
rect 2372 2148 2376 2204
rect 2376 2148 2432 2204
rect 2432 2148 2436 2204
rect 2372 2144 2436 2148
rect 2452 2204 2516 2208
rect 2452 2148 2456 2204
rect 2456 2148 2512 2204
rect 2512 2148 2516 2204
rect 2452 2144 2516 2148
rect 6212 2204 6276 2208
rect 6212 2148 6216 2204
rect 6216 2148 6272 2204
rect 6272 2148 6276 2204
rect 6212 2144 6276 2148
rect 6292 2204 6356 2208
rect 6292 2148 6296 2204
rect 6296 2148 6352 2204
rect 6352 2148 6356 2204
rect 6292 2144 6356 2148
rect 6372 2204 6436 2208
rect 6372 2148 6376 2204
rect 6376 2148 6432 2204
rect 6432 2148 6436 2204
rect 6372 2144 6436 2148
rect 6452 2204 6516 2208
rect 6452 2148 6456 2204
rect 6456 2148 6512 2204
rect 6512 2148 6516 2204
rect 6452 2144 6516 2148
rect 10212 2204 10276 2208
rect 10212 2148 10216 2204
rect 10216 2148 10272 2204
rect 10272 2148 10276 2204
rect 10212 2144 10276 2148
rect 10292 2204 10356 2208
rect 10292 2148 10296 2204
rect 10296 2148 10352 2204
rect 10352 2148 10356 2204
rect 10292 2144 10356 2148
rect 10372 2204 10436 2208
rect 10372 2148 10376 2204
rect 10376 2148 10432 2204
rect 10432 2148 10436 2204
rect 10372 2144 10436 2148
rect 10452 2204 10516 2208
rect 10452 2148 10456 2204
rect 10456 2148 10512 2204
rect 10512 2148 10516 2204
rect 10452 2144 10516 2148
rect 14212 2204 14276 2208
rect 14212 2148 14216 2204
rect 14216 2148 14272 2204
rect 14272 2148 14276 2204
rect 14212 2144 14276 2148
rect 14292 2204 14356 2208
rect 14292 2148 14296 2204
rect 14296 2148 14352 2204
rect 14352 2148 14356 2204
rect 14292 2144 14356 2148
rect 14372 2204 14436 2208
rect 14372 2148 14376 2204
rect 14376 2148 14432 2204
rect 14432 2148 14436 2204
rect 14372 2144 14436 2148
rect 14452 2204 14516 2208
rect 14452 2148 14456 2204
rect 14456 2148 14512 2204
rect 14512 2148 14516 2204
rect 14452 2144 14516 2148
rect 18212 2204 18276 2208
rect 18212 2148 18216 2204
rect 18216 2148 18272 2204
rect 18272 2148 18276 2204
rect 18212 2144 18276 2148
rect 18292 2204 18356 2208
rect 18292 2148 18296 2204
rect 18296 2148 18352 2204
rect 18352 2148 18356 2204
rect 18292 2144 18356 2148
rect 18372 2204 18436 2208
rect 18372 2148 18376 2204
rect 18376 2148 18432 2204
rect 18432 2148 18436 2204
rect 18372 2144 18436 2148
rect 18452 2204 18516 2208
rect 18452 2148 18456 2204
rect 18456 2148 18512 2204
rect 18512 2148 18516 2204
rect 18452 2144 18516 2148
<< metal4 >>
rect 1544 16896 1864 17456
rect 1544 16832 1552 16896
rect 1616 16832 1632 16896
rect 1696 16832 1712 16896
rect 1776 16832 1792 16896
rect 1856 16832 1864 16896
rect 1544 15808 1864 16832
rect 1544 15744 1552 15808
rect 1616 15744 1632 15808
rect 1696 15744 1712 15808
rect 1776 15744 1792 15808
rect 1856 15744 1864 15808
rect 1544 14894 1864 15744
rect 1544 14720 1586 14894
rect 1822 14720 1864 14894
rect 1544 14656 1552 14720
rect 1616 14656 1632 14658
rect 1696 14656 1712 14658
rect 1776 14656 1792 14658
rect 1856 14656 1864 14720
rect 1544 13632 1864 14656
rect 1544 13568 1552 13632
rect 1616 13568 1632 13632
rect 1696 13568 1712 13632
rect 1776 13568 1792 13632
rect 1856 13568 1864 13632
rect 1544 12544 1864 13568
rect 1544 12480 1552 12544
rect 1616 12480 1632 12544
rect 1696 12480 1712 12544
rect 1776 12480 1792 12544
rect 1856 12480 1864 12544
rect 1544 11456 1864 12480
rect 1544 11392 1552 11456
rect 1616 11392 1632 11456
rect 1696 11392 1712 11456
rect 1776 11392 1792 11456
rect 1856 11392 1864 11456
rect 1544 10894 1864 11392
rect 1544 10658 1586 10894
rect 1822 10658 1864 10894
rect 1544 10368 1864 10658
rect 1544 10304 1552 10368
rect 1616 10304 1632 10368
rect 1696 10304 1712 10368
rect 1776 10304 1792 10368
rect 1856 10304 1864 10368
rect 1544 9280 1864 10304
rect 1544 9216 1552 9280
rect 1616 9216 1632 9280
rect 1696 9216 1712 9280
rect 1776 9216 1792 9280
rect 1856 9216 1864 9280
rect 1544 8192 1864 9216
rect 1544 8128 1552 8192
rect 1616 8128 1632 8192
rect 1696 8128 1712 8192
rect 1776 8128 1792 8192
rect 1856 8128 1864 8192
rect 1544 7104 1864 8128
rect 1544 7040 1552 7104
rect 1616 7040 1632 7104
rect 1696 7040 1712 7104
rect 1776 7040 1792 7104
rect 1856 7040 1864 7104
rect 1544 6894 1864 7040
rect 1544 6658 1586 6894
rect 1822 6658 1864 6894
rect 1544 6016 1864 6658
rect 1544 5952 1552 6016
rect 1616 5952 1632 6016
rect 1696 5952 1712 6016
rect 1776 5952 1792 6016
rect 1856 5952 1864 6016
rect 1544 4928 1864 5952
rect 1544 4864 1552 4928
rect 1616 4864 1632 4928
rect 1696 4864 1712 4928
rect 1776 4864 1792 4928
rect 1856 4864 1864 4928
rect 1544 3840 1864 4864
rect 1544 3776 1552 3840
rect 1616 3776 1632 3840
rect 1696 3776 1712 3840
rect 1776 3776 1792 3840
rect 1856 3776 1864 3840
rect 1544 2894 1864 3776
rect 1544 2752 1586 2894
rect 1822 2752 1864 2894
rect 1544 2688 1552 2752
rect 1856 2688 1864 2752
rect 1544 2658 1586 2688
rect 1822 2658 1864 2688
rect 1544 2128 1864 2658
rect 2204 17440 2524 17456
rect 2204 17376 2212 17440
rect 2276 17376 2292 17440
rect 2356 17376 2372 17440
rect 2436 17376 2452 17440
rect 2516 17376 2524 17440
rect 2204 16352 2524 17376
rect 2204 16288 2212 16352
rect 2276 16288 2292 16352
rect 2356 16288 2372 16352
rect 2436 16288 2452 16352
rect 2516 16288 2524 16352
rect 2204 15554 2524 16288
rect 2204 15318 2246 15554
rect 2482 15318 2524 15554
rect 2204 15264 2524 15318
rect 2204 15200 2212 15264
rect 2276 15200 2292 15264
rect 2356 15200 2372 15264
rect 2436 15200 2452 15264
rect 2516 15200 2524 15264
rect 2204 14176 2524 15200
rect 2204 14112 2212 14176
rect 2276 14112 2292 14176
rect 2356 14112 2372 14176
rect 2436 14112 2452 14176
rect 2516 14112 2524 14176
rect 2204 13088 2524 14112
rect 2204 13024 2212 13088
rect 2276 13024 2292 13088
rect 2356 13024 2372 13088
rect 2436 13024 2452 13088
rect 2516 13024 2524 13088
rect 2204 12000 2524 13024
rect 2204 11936 2212 12000
rect 2276 11936 2292 12000
rect 2356 11936 2372 12000
rect 2436 11936 2452 12000
rect 2516 11936 2524 12000
rect 2204 11554 2524 11936
rect 2204 11318 2246 11554
rect 2482 11318 2524 11554
rect 2204 10912 2524 11318
rect 2204 10848 2212 10912
rect 2276 10848 2292 10912
rect 2356 10848 2372 10912
rect 2436 10848 2452 10912
rect 2516 10848 2524 10912
rect 2204 9824 2524 10848
rect 2204 9760 2212 9824
rect 2276 9760 2292 9824
rect 2356 9760 2372 9824
rect 2436 9760 2452 9824
rect 2516 9760 2524 9824
rect 2204 8736 2524 9760
rect 2204 8672 2212 8736
rect 2276 8672 2292 8736
rect 2356 8672 2372 8736
rect 2436 8672 2452 8736
rect 2516 8672 2524 8736
rect 2204 7648 2524 8672
rect 2204 7584 2212 7648
rect 2276 7584 2292 7648
rect 2356 7584 2372 7648
rect 2436 7584 2452 7648
rect 2516 7584 2524 7648
rect 2204 7554 2524 7584
rect 2204 7318 2246 7554
rect 2482 7318 2524 7554
rect 2204 6560 2524 7318
rect 2204 6496 2212 6560
rect 2276 6496 2292 6560
rect 2356 6496 2372 6560
rect 2436 6496 2452 6560
rect 2516 6496 2524 6560
rect 2204 5472 2524 6496
rect 2204 5408 2212 5472
rect 2276 5408 2292 5472
rect 2356 5408 2372 5472
rect 2436 5408 2452 5472
rect 2516 5408 2524 5472
rect 2204 4384 2524 5408
rect 2204 4320 2212 4384
rect 2276 4320 2292 4384
rect 2356 4320 2372 4384
rect 2436 4320 2452 4384
rect 2516 4320 2524 4384
rect 2204 3554 2524 4320
rect 2204 3318 2246 3554
rect 2482 3318 2524 3554
rect 2204 3296 2524 3318
rect 2204 3232 2212 3296
rect 2276 3232 2292 3296
rect 2356 3232 2372 3296
rect 2436 3232 2452 3296
rect 2516 3232 2524 3296
rect 2204 2208 2524 3232
rect 2204 2144 2212 2208
rect 2276 2144 2292 2208
rect 2356 2144 2372 2208
rect 2436 2144 2452 2208
rect 2516 2144 2524 2208
rect 2204 2128 2524 2144
rect 5544 16896 5864 17456
rect 5544 16832 5552 16896
rect 5616 16832 5632 16896
rect 5696 16832 5712 16896
rect 5776 16832 5792 16896
rect 5856 16832 5864 16896
rect 5544 15808 5864 16832
rect 5544 15744 5552 15808
rect 5616 15744 5632 15808
rect 5696 15744 5712 15808
rect 5776 15744 5792 15808
rect 5856 15744 5864 15808
rect 5544 14894 5864 15744
rect 5544 14720 5586 14894
rect 5822 14720 5864 14894
rect 5544 14656 5552 14720
rect 5616 14656 5632 14658
rect 5696 14656 5712 14658
rect 5776 14656 5792 14658
rect 5856 14656 5864 14720
rect 5544 13632 5864 14656
rect 5544 13568 5552 13632
rect 5616 13568 5632 13632
rect 5696 13568 5712 13632
rect 5776 13568 5792 13632
rect 5856 13568 5864 13632
rect 5544 12544 5864 13568
rect 5544 12480 5552 12544
rect 5616 12480 5632 12544
rect 5696 12480 5712 12544
rect 5776 12480 5792 12544
rect 5856 12480 5864 12544
rect 5544 11456 5864 12480
rect 5544 11392 5552 11456
rect 5616 11392 5632 11456
rect 5696 11392 5712 11456
rect 5776 11392 5792 11456
rect 5856 11392 5864 11456
rect 5544 10894 5864 11392
rect 5544 10658 5586 10894
rect 5822 10658 5864 10894
rect 5544 10368 5864 10658
rect 5544 10304 5552 10368
rect 5616 10304 5632 10368
rect 5696 10304 5712 10368
rect 5776 10304 5792 10368
rect 5856 10304 5864 10368
rect 5544 9280 5864 10304
rect 5544 9216 5552 9280
rect 5616 9216 5632 9280
rect 5696 9216 5712 9280
rect 5776 9216 5792 9280
rect 5856 9216 5864 9280
rect 5544 8192 5864 9216
rect 5544 8128 5552 8192
rect 5616 8128 5632 8192
rect 5696 8128 5712 8192
rect 5776 8128 5792 8192
rect 5856 8128 5864 8192
rect 5544 7104 5864 8128
rect 5544 7040 5552 7104
rect 5616 7040 5632 7104
rect 5696 7040 5712 7104
rect 5776 7040 5792 7104
rect 5856 7040 5864 7104
rect 5544 6894 5864 7040
rect 5544 6658 5586 6894
rect 5822 6658 5864 6894
rect 5544 6016 5864 6658
rect 5544 5952 5552 6016
rect 5616 5952 5632 6016
rect 5696 5952 5712 6016
rect 5776 5952 5792 6016
rect 5856 5952 5864 6016
rect 5544 4928 5864 5952
rect 5544 4864 5552 4928
rect 5616 4864 5632 4928
rect 5696 4864 5712 4928
rect 5776 4864 5792 4928
rect 5856 4864 5864 4928
rect 5544 3840 5864 4864
rect 5544 3776 5552 3840
rect 5616 3776 5632 3840
rect 5696 3776 5712 3840
rect 5776 3776 5792 3840
rect 5856 3776 5864 3840
rect 5544 2894 5864 3776
rect 5544 2752 5586 2894
rect 5822 2752 5864 2894
rect 5544 2688 5552 2752
rect 5856 2688 5864 2752
rect 5544 2658 5586 2688
rect 5822 2658 5864 2688
rect 5544 2128 5864 2658
rect 6204 17440 6524 17456
rect 6204 17376 6212 17440
rect 6276 17376 6292 17440
rect 6356 17376 6372 17440
rect 6436 17376 6452 17440
rect 6516 17376 6524 17440
rect 6204 16352 6524 17376
rect 6204 16288 6212 16352
rect 6276 16288 6292 16352
rect 6356 16288 6372 16352
rect 6436 16288 6452 16352
rect 6516 16288 6524 16352
rect 6204 15554 6524 16288
rect 6204 15318 6246 15554
rect 6482 15318 6524 15554
rect 6204 15264 6524 15318
rect 6204 15200 6212 15264
rect 6276 15200 6292 15264
rect 6356 15200 6372 15264
rect 6436 15200 6452 15264
rect 6516 15200 6524 15264
rect 6204 14176 6524 15200
rect 6204 14112 6212 14176
rect 6276 14112 6292 14176
rect 6356 14112 6372 14176
rect 6436 14112 6452 14176
rect 6516 14112 6524 14176
rect 6204 13088 6524 14112
rect 6204 13024 6212 13088
rect 6276 13024 6292 13088
rect 6356 13024 6372 13088
rect 6436 13024 6452 13088
rect 6516 13024 6524 13088
rect 6204 12000 6524 13024
rect 6204 11936 6212 12000
rect 6276 11936 6292 12000
rect 6356 11936 6372 12000
rect 6436 11936 6452 12000
rect 6516 11936 6524 12000
rect 6204 11554 6524 11936
rect 6204 11318 6246 11554
rect 6482 11318 6524 11554
rect 6204 10912 6524 11318
rect 6204 10848 6212 10912
rect 6276 10848 6292 10912
rect 6356 10848 6372 10912
rect 6436 10848 6452 10912
rect 6516 10848 6524 10912
rect 6204 9824 6524 10848
rect 6204 9760 6212 9824
rect 6276 9760 6292 9824
rect 6356 9760 6372 9824
rect 6436 9760 6452 9824
rect 6516 9760 6524 9824
rect 6204 8736 6524 9760
rect 6204 8672 6212 8736
rect 6276 8672 6292 8736
rect 6356 8672 6372 8736
rect 6436 8672 6452 8736
rect 6516 8672 6524 8736
rect 6204 7648 6524 8672
rect 6204 7584 6212 7648
rect 6276 7584 6292 7648
rect 6356 7584 6372 7648
rect 6436 7584 6452 7648
rect 6516 7584 6524 7648
rect 6204 7554 6524 7584
rect 6204 7318 6246 7554
rect 6482 7318 6524 7554
rect 6204 6560 6524 7318
rect 6204 6496 6212 6560
rect 6276 6496 6292 6560
rect 6356 6496 6372 6560
rect 6436 6496 6452 6560
rect 6516 6496 6524 6560
rect 6204 5472 6524 6496
rect 6204 5408 6212 5472
rect 6276 5408 6292 5472
rect 6356 5408 6372 5472
rect 6436 5408 6452 5472
rect 6516 5408 6524 5472
rect 6204 4384 6524 5408
rect 6204 4320 6212 4384
rect 6276 4320 6292 4384
rect 6356 4320 6372 4384
rect 6436 4320 6452 4384
rect 6516 4320 6524 4384
rect 6204 3554 6524 4320
rect 6204 3318 6246 3554
rect 6482 3318 6524 3554
rect 6204 3296 6524 3318
rect 6204 3232 6212 3296
rect 6276 3232 6292 3296
rect 6356 3232 6372 3296
rect 6436 3232 6452 3296
rect 6516 3232 6524 3296
rect 6204 2208 6524 3232
rect 6204 2144 6212 2208
rect 6276 2144 6292 2208
rect 6356 2144 6372 2208
rect 6436 2144 6452 2208
rect 6516 2144 6524 2208
rect 6204 2128 6524 2144
rect 9544 16896 9864 17456
rect 9544 16832 9552 16896
rect 9616 16832 9632 16896
rect 9696 16832 9712 16896
rect 9776 16832 9792 16896
rect 9856 16832 9864 16896
rect 9544 15808 9864 16832
rect 9544 15744 9552 15808
rect 9616 15744 9632 15808
rect 9696 15744 9712 15808
rect 9776 15744 9792 15808
rect 9856 15744 9864 15808
rect 9544 14894 9864 15744
rect 9544 14720 9586 14894
rect 9822 14720 9864 14894
rect 9544 14656 9552 14720
rect 9616 14656 9632 14658
rect 9696 14656 9712 14658
rect 9776 14656 9792 14658
rect 9856 14656 9864 14720
rect 9544 13632 9864 14656
rect 9544 13568 9552 13632
rect 9616 13568 9632 13632
rect 9696 13568 9712 13632
rect 9776 13568 9792 13632
rect 9856 13568 9864 13632
rect 9544 12544 9864 13568
rect 9544 12480 9552 12544
rect 9616 12480 9632 12544
rect 9696 12480 9712 12544
rect 9776 12480 9792 12544
rect 9856 12480 9864 12544
rect 9544 11456 9864 12480
rect 9544 11392 9552 11456
rect 9616 11392 9632 11456
rect 9696 11392 9712 11456
rect 9776 11392 9792 11456
rect 9856 11392 9864 11456
rect 9544 10894 9864 11392
rect 9544 10658 9586 10894
rect 9822 10658 9864 10894
rect 9544 10368 9864 10658
rect 9544 10304 9552 10368
rect 9616 10304 9632 10368
rect 9696 10304 9712 10368
rect 9776 10304 9792 10368
rect 9856 10304 9864 10368
rect 9544 9280 9864 10304
rect 9544 9216 9552 9280
rect 9616 9216 9632 9280
rect 9696 9216 9712 9280
rect 9776 9216 9792 9280
rect 9856 9216 9864 9280
rect 9544 8192 9864 9216
rect 9544 8128 9552 8192
rect 9616 8128 9632 8192
rect 9696 8128 9712 8192
rect 9776 8128 9792 8192
rect 9856 8128 9864 8192
rect 9544 7104 9864 8128
rect 9544 7040 9552 7104
rect 9616 7040 9632 7104
rect 9696 7040 9712 7104
rect 9776 7040 9792 7104
rect 9856 7040 9864 7104
rect 9544 6894 9864 7040
rect 9544 6658 9586 6894
rect 9822 6658 9864 6894
rect 9544 6016 9864 6658
rect 9544 5952 9552 6016
rect 9616 5952 9632 6016
rect 9696 5952 9712 6016
rect 9776 5952 9792 6016
rect 9856 5952 9864 6016
rect 9544 4928 9864 5952
rect 9544 4864 9552 4928
rect 9616 4864 9632 4928
rect 9696 4864 9712 4928
rect 9776 4864 9792 4928
rect 9856 4864 9864 4928
rect 9544 3840 9864 4864
rect 9544 3776 9552 3840
rect 9616 3776 9632 3840
rect 9696 3776 9712 3840
rect 9776 3776 9792 3840
rect 9856 3776 9864 3840
rect 9544 2894 9864 3776
rect 9544 2752 9586 2894
rect 9822 2752 9864 2894
rect 9544 2688 9552 2752
rect 9856 2688 9864 2752
rect 9544 2658 9586 2688
rect 9822 2658 9864 2688
rect 9544 2128 9864 2658
rect 10204 17440 10524 17456
rect 10204 17376 10212 17440
rect 10276 17376 10292 17440
rect 10356 17376 10372 17440
rect 10436 17376 10452 17440
rect 10516 17376 10524 17440
rect 10204 16352 10524 17376
rect 10204 16288 10212 16352
rect 10276 16288 10292 16352
rect 10356 16288 10372 16352
rect 10436 16288 10452 16352
rect 10516 16288 10524 16352
rect 10204 15554 10524 16288
rect 10204 15318 10246 15554
rect 10482 15318 10524 15554
rect 10204 15264 10524 15318
rect 10204 15200 10212 15264
rect 10276 15200 10292 15264
rect 10356 15200 10372 15264
rect 10436 15200 10452 15264
rect 10516 15200 10524 15264
rect 10204 14176 10524 15200
rect 10204 14112 10212 14176
rect 10276 14112 10292 14176
rect 10356 14112 10372 14176
rect 10436 14112 10452 14176
rect 10516 14112 10524 14176
rect 10204 13088 10524 14112
rect 10204 13024 10212 13088
rect 10276 13024 10292 13088
rect 10356 13024 10372 13088
rect 10436 13024 10452 13088
rect 10516 13024 10524 13088
rect 10204 12000 10524 13024
rect 10204 11936 10212 12000
rect 10276 11936 10292 12000
rect 10356 11936 10372 12000
rect 10436 11936 10452 12000
rect 10516 11936 10524 12000
rect 10204 11554 10524 11936
rect 10204 11318 10246 11554
rect 10482 11318 10524 11554
rect 10204 10912 10524 11318
rect 10204 10848 10212 10912
rect 10276 10848 10292 10912
rect 10356 10848 10372 10912
rect 10436 10848 10452 10912
rect 10516 10848 10524 10912
rect 10204 9824 10524 10848
rect 10204 9760 10212 9824
rect 10276 9760 10292 9824
rect 10356 9760 10372 9824
rect 10436 9760 10452 9824
rect 10516 9760 10524 9824
rect 10204 8736 10524 9760
rect 10204 8672 10212 8736
rect 10276 8672 10292 8736
rect 10356 8672 10372 8736
rect 10436 8672 10452 8736
rect 10516 8672 10524 8736
rect 10204 7648 10524 8672
rect 10204 7584 10212 7648
rect 10276 7584 10292 7648
rect 10356 7584 10372 7648
rect 10436 7584 10452 7648
rect 10516 7584 10524 7648
rect 10204 7554 10524 7584
rect 10204 7318 10246 7554
rect 10482 7318 10524 7554
rect 10204 6560 10524 7318
rect 10204 6496 10212 6560
rect 10276 6496 10292 6560
rect 10356 6496 10372 6560
rect 10436 6496 10452 6560
rect 10516 6496 10524 6560
rect 10204 5472 10524 6496
rect 10204 5408 10212 5472
rect 10276 5408 10292 5472
rect 10356 5408 10372 5472
rect 10436 5408 10452 5472
rect 10516 5408 10524 5472
rect 10204 4384 10524 5408
rect 10204 4320 10212 4384
rect 10276 4320 10292 4384
rect 10356 4320 10372 4384
rect 10436 4320 10452 4384
rect 10516 4320 10524 4384
rect 10204 3554 10524 4320
rect 10204 3318 10246 3554
rect 10482 3318 10524 3554
rect 10204 3296 10524 3318
rect 10204 3232 10212 3296
rect 10276 3232 10292 3296
rect 10356 3232 10372 3296
rect 10436 3232 10452 3296
rect 10516 3232 10524 3296
rect 10204 2208 10524 3232
rect 10204 2144 10212 2208
rect 10276 2144 10292 2208
rect 10356 2144 10372 2208
rect 10436 2144 10452 2208
rect 10516 2144 10524 2208
rect 10204 2128 10524 2144
rect 13544 16896 13864 17456
rect 13544 16832 13552 16896
rect 13616 16832 13632 16896
rect 13696 16832 13712 16896
rect 13776 16832 13792 16896
rect 13856 16832 13864 16896
rect 13544 15808 13864 16832
rect 13544 15744 13552 15808
rect 13616 15744 13632 15808
rect 13696 15744 13712 15808
rect 13776 15744 13792 15808
rect 13856 15744 13864 15808
rect 13544 14894 13864 15744
rect 13544 14720 13586 14894
rect 13822 14720 13864 14894
rect 13544 14656 13552 14720
rect 13616 14656 13632 14658
rect 13696 14656 13712 14658
rect 13776 14656 13792 14658
rect 13856 14656 13864 14720
rect 13544 13632 13864 14656
rect 13544 13568 13552 13632
rect 13616 13568 13632 13632
rect 13696 13568 13712 13632
rect 13776 13568 13792 13632
rect 13856 13568 13864 13632
rect 13544 12544 13864 13568
rect 13544 12480 13552 12544
rect 13616 12480 13632 12544
rect 13696 12480 13712 12544
rect 13776 12480 13792 12544
rect 13856 12480 13864 12544
rect 13544 11456 13864 12480
rect 13544 11392 13552 11456
rect 13616 11392 13632 11456
rect 13696 11392 13712 11456
rect 13776 11392 13792 11456
rect 13856 11392 13864 11456
rect 13544 10894 13864 11392
rect 13544 10658 13586 10894
rect 13822 10658 13864 10894
rect 13544 10368 13864 10658
rect 13544 10304 13552 10368
rect 13616 10304 13632 10368
rect 13696 10304 13712 10368
rect 13776 10304 13792 10368
rect 13856 10304 13864 10368
rect 13544 9280 13864 10304
rect 13544 9216 13552 9280
rect 13616 9216 13632 9280
rect 13696 9216 13712 9280
rect 13776 9216 13792 9280
rect 13856 9216 13864 9280
rect 13544 8192 13864 9216
rect 13544 8128 13552 8192
rect 13616 8128 13632 8192
rect 13696 8128 13712 8192
rect 13776 8128 13792 8192
rect 13856 8128 13864 8192
rect 13544 7104 13864 8128
rect 13544 7040 13552 7104
rect 13616 7040 13632 7104
rect 13696 7040 13712 7104
rect 13776 7040 13792 7104
rect 13856 7040 13864 7104
rect 13544 6894 13864 7040
rect 13544 6658 13586 6894
rect 13822 6658 13864 6894
rect 13544 6016 13864 6658
rect 13544 5952 13552 6016
rect 13616 5952 13632 6016
rect 13696 5952 13712 6016
rect 13776 5952 13792 6016
rect 13856 5952 13864 6016
rect 13544 4928 13864 5952
rect 13544 4864 13552 4928
rect 13616 4864 13632 4928
rect 13696 4864 13712 4928
rect 13776 4864 13792 4928
rect 13856 4864 13864 4928
rect 13544 3840 13864 4864
rect 13544 3776 13552 3840
rect 13616 3776 13632 3840
rect 13696 3776 13712 3840
rect 13776 3776 13792 3840
rect 13856 3776 13864 3840
rect 13544 2894 13864 3776
rect 13544 2752 13586 2894
rect 13822 2752 13864 2894
rect 13544 2688 13552 2752
rect 13856 2688 13864 2752
rect 13544 2658 13586 2688
rect 13822 2658 13864 2688
rect 13544 2128 13864 2658
rect 14204 17440 14524 17456
rect 14204 17376 14212 17440
rect 14276 17376 14292 17440
rect 14356 17376 14372 17440
rect 14436 17376 14452 17440
rect 14516 17376 14524 17440
rect 14204 16352 14524 17376
rect 14204 16288 14212 16352
rect 14276 16288 14292 16352
rect 14356 16288 14372 16352
rect 14436 16288 14452 16352
rect 14516 16288 14524 16352
rect 14204 15554 14524 16288
rect 14204 15318 14246 15554
rect 14482 15318 14524 15554
rect 14204 15264 14524 15318
rect 14204 15200 14212 15264
rect 14276 15200 14292 15264
rect 14356 15200 14372 15264
rect 14436 15200 14452 15264
rect 14516 15200 14524 15264
rect 14204 14176 14524 15200
rect 14204 14112 14212 14176
rect 14276 14112 14292 14176
rect 14356 14112 14372 14176
rect 14436 14112 14452 14176
rect 14516 14112 14524 14176
rect 14204 13088 14524 14112
rect 14204 13024 14212 13088
rect 14276 13024 14292 13088
rect 14356 13024 14372 13088
rect 14436 13024 14452 13088
rect 14516 13024 14524 13088
rect 14204 12000 14524 13024
rect 14204 11936 14212 12000
rect 14276 11936 14292 12000
rect 14356 11936 14372 12000
rect 14436 11936 14452 12000
rect 14516 11936 14524 12000
rect 14204 11554 14524 11936
rect 14204 11318 14246 11554
rect 14482 11318 14524 11554
rect 14204 10912 14524 11318
rect 14204 10848 14212 10912
rect 14276 10848 14292 10912
rect 14356 10848 14372 10912
rect 14436 10848 14452 10912
rect 14516 10848 14524 10912
rect 14204 9824 14524 10848
rect 14204 9760 14212 9824
rect 14276 9760 14292 9824
rect 14356 9760 14372 9824
rect 14436 9760 14452 9824
rect 14516 9760 14524 9824
rect 14204 8736 14524 9760
rect 14204 8672 14212 8736
rect 14276 8672 14292 8736
rect 14356 8672 14372 8736
rect 14436 8672 14452 8736
rect 14516 8672 14524 8736
rect 14204 7648 14524 8672
rect 14204 7584 14212 7648
rect 14276 7584 14292 7648
rect 14356 7584 14372 7648
rect 14436 7584 14452 7648
rect 14516 7584 14524 7648
rect 14204 7554 14524 7584
rect 14204 7318 14246 7554
rect 14482 7318 14524 7554
rect 14204 6560 14524 7318
rect 14204 6496 14212 6560
rect 14276 6496 14292 6560
rect 14356 6496 14372 6560
rect 14436 6496 14452 6560
rect 14516 6496 14524 6560
rect 14204 5472 14524 6496
rect 14204 5408 14212 5472
rect 14276 5408 14292 5472
rect 14356 5408 14372 5472
rect 14436 5408 14452 5472
rect 14516 5408 14524 5472
rect 14204 4384 14524 5408
rect 14204 4320 14212 4384
rect 14276 4320 14292 4384
rect 14356 4320 14372 4384
rect 14436 4320 14452 4384
rect 14516 4320 14524 4384
rect 14204 3554 14524 4320
rect 14204 3318 14246 3554
rect 14482 3318 14524 3554
rect 14204 3296 14524 3318
rect 14204 3232 14212 3296
rect 14276 3232 14292 3296
rect 14356 3232 14372 3296
rect 14436 3232 14452 3296
rect 14516 3232 14524 3296
rect 14204 2208 14524 3232
rect 14204 2144 14212 2208
rect 14276 2144 14292 2208
rect 14356 2144 14372 2208
rect 14436 2144 14452 2208
rect 14516 2144 14524 2208
rect 14204 2128 14524 2144
rect 17544 16896 17864 17456
rect 17544 16832 17552 16896
rect 17616 16832 17632 16896
rect 17696 16832 17712 16896
rect 17776 16832 17792 16896
rect 17856 16832 17864 16896
rect 17544 15808 17864 16832
rect 17544 15744 17552 15808
rect 17616 15744 17632 15808
rect 17696 15744 17712 15808
rect 17776 15744 17792 15808
rect 17856 15744 17864 15808
rect 17544 14894 17864 15744
rect 17544 14720 17586 14894
rect 17822 14720 17864 14894
rect 17544 14656 17552 14720
rect 17616 14656 17632 14658
rect 17696 14656 17712 14658
rect 17776 14656 17792 14658
rect 17856 14656 17864 14720
rect 17544 13632 17864 14656
rect 17544 13568 17552 13632
rect 17616 13568 17632 13632
rect 17696 13568 17712 13632
rect 17776 13568 17792 13632
rect 17856 13568 17864 13632
rect 17544 12544 17864 13568
rect 17544 12480 17552 12544
rect 17616 12480 17632 12544
rect 17696 12480 17712 12544
rect 17776 12480 17792 12544
rect 17856 12480 17864 12544
rect 17544 11456 17864 12480
rect 17544 11392 17552 11456
rect 17616 11392 17632 11456
rect 17696 11392 17712 11456
rect 17776 11392 17792 11456
rect 17856 11392 17864 11456
rect 17544 10894 17864 11392
rect 17544 10658 17586 10894
rect 17822 10658 17864 10894
rect 17544 10368 17864 10658
rect 17544 10304 17552 10368
rect 17616 10304 17632 10368
rect 17696 10304 17712 10368
rect 17776 10304 17792 10368
rect 17856 10304 17864 10368
rect 17544 9280 17864 10304
rect 17544 9216 17552 9280
rect 17616 9216 17632 9280
rect 17696 9216 17712 9280
rect 17776 9216 17792 9280
rect 17856 9216 17864 9280
rect 17544 8192 17864 9216
rect 17544 8128 17552 8192
rect 17616 8128 17632 8192
rect 17696 8128 17712 8192
rect 17776 8128 17792 8192
rect 17856 8128 17864 8192
rect 17544 7104 17864 8128
rect 17544 7040 17552 7104
rect 17616 7040 17632 7104
rect 17696 7040 17712 7104
rect 17776 7040 17792 7104
rect 17856 7040 17864 7104
rect 17544 6894 17864 7040
rect 17544 6658 17586 6894
rect 17822 6658 17864 6894
rect 17544 6016 17864 6658
rect 17544 5952 17552 6016
rect 17616 5952 17632 6016
rect 17696 5952 17712 6016
rect 17776 5952 17792 6016
rect 17856 5952 17864 6016
rect 17544 4928 17864 5952
rect 17544 4864 17552 4928
rect 17616 4864 17632 4928
rect 17696 4864 17712 4928
rect 17776 4864 17792 4928
rect 17856 4864 17864 4928
rect 17544 3840 17864 4864
rect 17544 3776 17552 3840
rect 17616 3776 17632 3840
rect 17696 3776 17712 3840
rect 17776 3776 17792 3840
rect 17856 3776 17864 3840
rect 17544 2894 17864 3776
rect 17544 2752 17586 2894
rect 17822 2752 17864 2894
rect 17544 2688 17552 2752
rect 17856 2688 17864 2752
rect 17544 2658 17586 2688
rect 17822 2658 17864 2688
rect 17544 2128 17864 2658
rect 18204 17440 18524 17456
rect 18204 17376 18212 17440
rect 18276 17376 18292 17440
rect 18356 17376 18372 17440
rect 18436 17376 18452 17440
rect 18516 17376 18524 17440
rect 18204 16352 18524 17376
rect 18204 16288 18212 16352
rect 18276 16288 18292 16352
rect 18356 16288 18372 16352
rect 18436 16288 18452 16352
rect 18516 16288 18524 16352
rect 18204 15554 18524 16288
rect 18204 15318 18246 15554
rect 18482 15318 18524 15554
rect 18204 15264 18524 15318
rect 18204 15200 18212 15264
rect 18276 15200 18292 15264
rect 18356 15200 18372 15264
rect 18436 15200 18452 15264
rect 18516 15200 18524 15264
rect 18204 14176 18524 15200
rect 18204 14112 18212 14176
rect 18276 14112 18292 14176
rect 18356 14112 18372 14176
rect 18436 14112 18452 14176
rect 18516 14112 18524 14176
rect 18204 13088 18524 14112
rect 18204 13024 18212 13088
rect 18276 13024 18292 13088
rect 18356 13024 18372 13088
rect 18436 13024 18452 13088
rect 18516 13024 18524 13088
rect 18204 12000 18524 13024
rect 18204 11936 18212 12000
rect 18276 11936 18292 12000
rect 18356 11936 18372 12000
rect 18436 11936 18452 12000
rect 18516 11936 18524 12000
rect 18204 11554 18524 11936
rect 18204 11318 18246 11554
rect 18482 11318 18524 11554
rect 18204 10912 18524 11318
rect 18204 10848 18212 10912
rect 18276 10848 18292 10912
rect 18356 10848 18372 10912
rect 18436 10848 18452 10912
rect 18516 10848 18524 10912
rect 18204 9824 18524 10848
rect 18204 9760 18212 9824
rect 18276 9760 18292 9824
rect 18356 9760 18372 9824
rect 18436 9760 18452 9824
rect 18516 9760 18524 9824
rect 18204 8736 18524 9760
rect 18204 8672 18212 8736
rect 18276 8672 18292 8736
rect 18356 8672 18372 8736
rect 18436 8672 18452 8736
rect 18516 8672 18524 8736
rect 18204 7648 18524 8672
rect 18204 7584 18212 7648
rect 18276 7584 18292 7648
rect 18356 7584 18372 7648
rect 18436 7584 18452 7648
rect 18516 7584 18524 7648
rect 18204 7554 18524 7584
rect 18204 7318 18246 7554
rect 18482 7318 18524 7554
rect 18204 6560 18524 7318
rect 18204 6496 18212 6560
rect 18276 6496 18292 6560
rect 18356 6496 18372 6560
rect 18436 6496 18452 6560
rect 18516 6496 18524 6560
rect 18204 5472 18524 6496
rect 18204 5408 18212 5472
rect 18276 5408 18292 5472
rect 18356 5408 18372 5472
rect 18436 5408 18452 5472
rect 18516 5408 18524 5472
rect 18204 4384 18524 5408
rect 18204 4320 18212 4384
rect 18276 4320 18292 4384
rect 18356 4320 18372 4384
rect 18436 4320 18452 4384
rect 18516 4320 18524 4384
rect 18204 3554 18524 4320
rect 18204 3318 18246 3554
rect 18482 3318 18524 3554
rect 18204 3296 18524 3318
rect 18204 3232 18212 3296
rect 18276 3232 18292 3296
rect 18356 3232 18372 3296
rect 18436 3232 18452 3296
rect 18516 3232 18524 3296
rect 18204 2208 18524 3232
rect 18204 2144 18212 2208
rect 18276 2144 18292 2208
rect 18356 2144 18372 2208
rect 18436 2144 18452 2208
rect 18516 2144 18524 2208
rect 18204 2128 18524 2144
<< via4 >>
rect 1586 14720 1822 14894
rect 1586 14658 1616 14720
rect 1616 14658 1632 14720
rect 1632 14658 1696 14720
rect 1696 14658 1712 14720
rect 1712 14658 1776 14720
rect 1776 14658 1792 14720
rect 1792 14658 1822 14720
rect 1586 10658 1822 10894
rect 1586 6658 1822 6894
rect 1586 2752 1822 2894
rect 1586 2688 1616 2752
rect 1616 2688 1632 2752
rect 1632 2688 1696 2752
rect 1696 2688 1712 2752
rect 1712 2688 1776 2752
rect 1776 2688 1792 2752
rect 1792 2688 1822 2752
rect 1586 2658 1822 2688
rect 2246 15318 2482 15554
rect 2246 11318 2482 11554
rect 2246 7318 2482 7554
rect 2246 3318 2482 3554
rect 5586 14720 5822 14894
rect 5586 14658 5616 14720
rect 5616 14658 5632 14720
rect 5632 14658 5696 14720
rect 5696 14658 5712 14720
rect 5712 14658 5776 14720
rect 5776 14658 5792 14720
rect 5792 14658 5822 14720
rect 5586 10658 5822 10894
rect 5586 6658 5822 6894
rect 5586 2752 5822 2894
rect 5586 2688 5616 2752
rect 5616 2688 5632 2752
rect 5632 2688 5696 2752
rect 5696 2688 5712 2752
rect 5712 2688 5776 2752
rect 5776 2688 5792 2752
rect 5792 2688 5822 2752
rect 5586 2658 5822 2688
rect 6246 15318 6482 15554
rect 6246 11318 6482 11554
rect 6246 7318 6482 7554
rect 6246 3318 6482 3554
rect 9586 14720 9822 14894
rect 9586 14658 9616 14720
rect 9616 14658 9632 14720
rect 9632 14658 9696 14720
rect 9696 14658 9712 14720
rect 9712 14658 9776 14720
rect 9776 14658 9792 14720
rect 9792 14658 9822 14720
rect 9586 10658 9822 10894
rect 9586 6658 9822 6894
rect 9586 2752 9822 2894
rect 9586 2688 9616 2752
rect 9616 2688 9632 2752
rect 9632 2688 9696 2752
rect 9696 2688 9712 2752
rect 9712 2688 9776 2752
rect 9776 2688 9792 2752
rect 9792 2688 9822 2752
rect 9586 2658 9822 2688
rect 10246 15318 10482 15554
rect 10246 11318 10482 11554
rect 10246 7318 10482 7554
rect 10246 3318 10482 3554
rect 13586 14720 13822 14894
rect 13586 14658 13616 14720
rect 13616 14658 13632 14720
rect 13632 14658 13696 14720
rect 13696 14658 13712 14720
rect 13712 14658 13776 14720
rect 13776 14658 13792 14720
rect 13792 14658 13822 14720
rect 13586 10658 13822 10894
rect 13586 6658 13822 6894
rect 13586 2752 13822 2894
rect 13586 2688 13616 2752
rect 13616 2688 13632 2752
rect 13632 2688 13696 2752
rect 13696 2688 13712 2752
rect 13712 2688 13776 2752
rect 13776 2688 13792 2752
rect 13792 2688 13822 2752
rect 13586 2658 13822 2688
rect 14246 15318 14482 15554
rect 14246 11318 14482 11554
rect 14246 7318 14482 7554
rect 14246 3318 14482 3554
rect 17586 14720 17822 14894
rect 17586 14658 17616 14720
rect 17616 14658 17632 14720
rect 17632 14658 17696 14720
rect 17696 14658 17712 14720
rect 17712 14658 17776 14720
rect 17776 14658 17792 14720
rect 17792 14658 17822 14720
rect 17586 10658 17822 10894
rect 17586 6658 17822 6894
rect 17586 2752 17822 2894
rect 17586 2688 17616 2752
rect 17616 2688 17632 2752
rect 17632 2688 17696 2752
rect 17696 2688 17712 2752
rect 17712 2688 17776 2752
rect 17776 2688 17792 2752
rect 17792 2688 17822 2752
rect 17586 2658 17822 2688
rect 18246 15318 18482 15554
rect 18246 11318 18482 11554
rect 18246 7318 18482 7554
rect 18246 3318 18482 3554
<< metal5 >>
rect 1056 15554 18908 15596
rect 1056 15318 2246 15554
rect 2482 15318 6246 15554
rect 6482 15318 10246 15554
rect 10482 15318 14246 15554
rect 14482 15318 18246 15554
rect 18482 15318 18908 15554
rect 1056 15276 18908 15318
rect 1056 14894 18908 14936
rect 1056 14658 1586 14894
rect 1822 14658 5586 14894
rect 5822 14658 9586 14894
rect 9822 14658 13586 14894
rect 13822 14658 17586 14894
rect 17822 14658 18908 14894
rect 1056 14616 18908 14658
rect 1056 11554 18908 11596
rect 1056 11318 2246 11554
rect 2482 11318 6246 11554
rect 6482 11318 10246 11554
rect 10482 11318 14246 11554
rect 14482 11318 18246 11554
rect 18482 11318 18908 11554
rect 1056 11276 18908 11318
rect 1056 10894 18908 10936
rect 1056 10658 1586 10894
rect 1822 10658 5586 10894
rect 5822 10658 9586 10894
rect 9822 10658 13586 10894
rect 13822 10658 17586 10894
rect 17822 10658 18908 10894
rect 1056 10616 18908 10658
rect 1056 7554 18908 7596
rect 1056 7318 2246 7554
rect 2482 7318 6246 7554
rect 6482 7318 10246 7554
rect 10482 7318 14246 7554
rect 14482 7318 18246 7554
rect 18482 7318 18908 7554
rect 1056 7276 18908 7318
rect 1056 6894 18908 6936
rect 1056 6658 1586 6894
rect 1822 6658 5586 6894
rect 5822 6658 9586 6894
rect 9822 6658 13586 6894
rect 13822 6658 17586 6894
rect 17822 6658 18908 6894
rect 1056 6616 18908 6658
rect 1056 3554 18908 3596
rect 1056 3318 2246 3554
rect 2482 3318 6246 3554
rect 6482 3318 10246 3554
rect 10482 3318 14246 3554
rect 14482 3318 18246 3554
rect 18482 3318 18908 3554
rect 1056 3276 18908 3318
rect 1056 2894 18908 2936
rect 1056 2658 1586 2894
rect 1822 2658 5586 2894
rect 5822 2658 9586 2894
rect 9822 2658 13586 2894
rect 13822 2658 17586 2894
rect 17822 2658 18908 2894
rect 1056 2616 18908 2658
use sky130_fd_sc_hd__conb_1  cpu_lab6_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_2
timestamp 1704896540
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_3
timestamp 1704896540
transform 1 0 18308 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_4
timestamp 1704896540
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_5
timestamp 1704896540
transform -1 0 10028 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_6
timestamp 1704896540
transform -1 0 10672 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_7
timestamp 1704896540
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_8
timestamp 1704896540
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_9
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_10
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  cpu_lab6_11
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1704896540
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_104
timestamp 1704896540
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_189
timestamp 1704896540
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1704896540
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 1704896540
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1704896540
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1704896540
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1704896540
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_189
timestamp 1704896540
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1704896540
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1704896540
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_181
timestamp 1704896540
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_189
timestamp 1704896540
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1704896540
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1704896540
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1704896540
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_189
timestamp 1704896540
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1704896540
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_189
timestamp 1704896540
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1704896540
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1704896540
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1704896540
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_189
timestamp 1704896540
transform 1 0 18492 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1704896540
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1704896540
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_181
timestamp 1704896540
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_189
timestamp 1704896540
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1704896540
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1704896540
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1704896540
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1704896540
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1704896540
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1704896540
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1704896540
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1704896540
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_189
timestamp 1704896540
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1704896540
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1704896540
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1704896540
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1704896540
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1704896540
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1704896540
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1704896540
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1704896540
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_181
timestamp 1704896540
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_189
timestamp 1704896540
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1704896540
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1704896540
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1704896540
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1704896540
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1704896540
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1704896540
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1704896540
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1704896540
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1704896540
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1704896540
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_189
timestamp 1704896540
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_6
timestamp 1704896540
transform 1 0 1656 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_18
timestamp 1704896540
transform 1 0 2760 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_30
timestamp 1704896540
transform 1 0 3864 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_42
timestamp 1704896540
transform 1 0 4968 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1704896540
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1704896540
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1704896540
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1704896540
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1704896540
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1704896540
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1704896540
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1704896540
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1704896540
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_181
timestamp 1704896540
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_189
timestamp 1704896540
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 1704896540
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 1704896540
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1704896540
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1704896540
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1704896540
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1704896540
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1704896540
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1704896540
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1704896540
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1704896540
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1704896540
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1704896540
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_189
timestamp 1704896540
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1704896540
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1704896540
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1704896540
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1704896540
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1704896540
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1704896540
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1704896540
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1704896540
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1704896540
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1704896540
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_181
timestamp 1704896540
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_189
timestamp 1704896540
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_6
timestamp 1704896540
transform 1 0 1656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_18
timestamp 1704896540
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1704896540
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1704896540
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1704896540
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1704896540
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1704896540
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1704896540
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1704896540
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1704896540
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1704896540
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1704896540
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1704896540
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1704896540
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_189
timestamp 1704896540
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_6
timestamp 1704896540
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_18
timestamp 1704896540
transform 1 0 2760 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_30
timestamp 1704896540
transform 1 0 3864 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_42
timestamp 1704896540
transform 1 0 4968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1704896540
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1704896540
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1704896540
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1704896540
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1704896540
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1704896540
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1704896540
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1704896540
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1704896540
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_181
timestamp 1704896540
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_6
timestamp 1704896540
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_18
timestamp 1704896540
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1704896540
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1704896540
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1704896540
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1704896540
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1704896540
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1704896540
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1704896540
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1704896540
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1704896540
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1704896540
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1704896540
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1704896540
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1704896540
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1704896540
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_189
timestamp 1704896540
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_6
timestamp 1704896540
transform 1 0 1656 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_18
timestamp 1704896540
transform 1 0 2760 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_30
timestamp 1704896540
transform 1 0 3864 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_42
timestamp 1704896540
transform 1 0 4968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1704896540
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1704896540
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1704896540
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1704896540
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1704896540
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1704896540
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1704896540
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1704896540
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1704896540
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1704896540
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1704896540
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1704896540
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1704896540
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_189
timestamp 1704896540
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1704896540
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1704896540
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1704896540
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1704896540
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1704896540
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1704896540
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1704896540
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1704896540
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1704896540
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1704896540
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1704896540
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1704896540
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_189
timestamp 1704896540
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1704896540
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1704896540
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1704896540
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1704896540
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1704896540
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1704896540
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1704896540
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1704896540
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1704896540
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1704896540
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1704896540
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1704896540
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1704896540
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1704896540
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_181
timestamp 1704896540
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_189
timestamp 1704896540
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1704896540
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1704896540
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1704896540
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1704896540
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1704896540
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1704896540
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1704896540
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1704896540
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1704896540
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1704896540
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1704896540
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_189
timestamp 1704896540
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1704896540
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1704896540
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1704896540
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1704896540
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1704896540
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1704896540
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1704896540
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1704896540
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1704896540
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1704896540
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1704896540
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1704896540
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1704896540
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_181
timestamp 1704896540
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 1704896540
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1704896540
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1704896540
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1704896540
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1704896540
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1704896540
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1704896540
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1704896540
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1704896540
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1704896540
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1704896540
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1704896540
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1704896540
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1704896540
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1704896540
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_189
timestamp 1704896540
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1704896540
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1704896540
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1704896540
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1704896540
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1704896540
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1704896540
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1704896540
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1704896540
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1704896540
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1704896540
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1704896540
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1704896540
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1704896540
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1704896540
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1704896540
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_181
timestamp 1704896540
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_189
timestamp 1704896540
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1704896540
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1704896540
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1704896540
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1704896540
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1704896540
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1704896540
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1704896540
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1704896540
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1704896540
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1704896540
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1704896540
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1704896540
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1704896540
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1704896540
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_189
timestamp 1704896540
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1704896540
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1704896540
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1704896540
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1704896540
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1704896540
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1704896540
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1704896540
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1704896540
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1704896540
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1704896540
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1704896540
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1704896540
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1704896540
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1704896540
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1704896540
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1704896540
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_181
timestamp 1704896540
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_189
timestamp 1704896540
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1704896540
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1704896540
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1704896540
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1704896540
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1704896540
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1704896540
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1704896540
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1704896540
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1704896540
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1704896540
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1704896540
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1704896540
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1704896540
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1704896540
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1704896540
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1704896540
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_189
timestamp 1704896540
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1704896540
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1704896540
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_27
timestamp 1704896540
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_29
timestamp 1704896540
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_41
timestamp 1704896540
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_53
timestamp 1704896540
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1704896540
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1704896540
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_81
timestamp 1704896540
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_85
timestamp 1704896540
transform 1 0 8924 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_93
timestamp 1704896540
transform 1 0 9660 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_97
timestamp 1704896540
transform 1 0 10028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_104
timestamp 1704896540
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1704896540
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1704896540
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_137
timestamp 1704896540
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_141
timestamp 1704896540
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_153
timestamp 1704896540
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1704896540
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_181
timestamp 1704896540
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_189
timestamp 1704896540
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_28
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_29
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_30
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_31
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_32
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_33
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_34
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_35
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_36
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_37
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_38
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_39
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_40
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_41
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_42
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_43
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_44
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_45
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_46
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_47
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_48
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_49
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_50
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_51
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_52
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_53
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_54
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_55
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_62
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_63
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_65
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_66
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_68
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_69
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_71
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_72
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_74
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_75
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_78
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_89
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_92
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_93
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_95
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_96
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_98
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_99
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_101
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_102
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_104
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_105
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_107
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_108
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_110
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_111
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_113
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_114
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_116
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_117
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_119
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_120
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_122
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_123
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_125
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_126
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_128
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_129
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_131
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_132
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_134
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_135
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_137
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_138
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_140
timestamp 1704896540
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_141
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 1704896540
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 1704896540
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_145
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
<< labels >>
flabel metal4 s 2204 2128 2524 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6204 2128 6524 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 10204 2128 10524 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 14204 2128 14524 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 18204 2128 18524 17456 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3276 18908 3596 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7276 18908 7596 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 11276 18908 11596 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 15276 18908 15596 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1544 2128 1864 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5544 2128 5864 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9544 2128 9864 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13544 2128 13864 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 17544 2128 17864 17456 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 2616 18908 2936 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 6616 18908 6936 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 10616 18908 10936 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 14616 18908 14936 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 an[0]
port 2 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 an[1]
port 3 nsew signal output
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 an[2]
port 4 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 an[3]
port 5 nsew signal output
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 clk
port 6 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 control
port 7 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 reset
port 8 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 seg[0]
port 9 nsew signal output
flabel metal3 s 19200 10208 20000 10328 0 FreeSans 480 0 0 0 seg[1]
port 10 nsew signal output
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 seg[2]
port 11 nsew signal output
flabel metal2 s 9678 19200 9734 20000 0 FreeSans 224 90 0 0 seg[3]
port 12 nsew signal output
flabel metal2 s 10322 19200 10378 20000 0 FreeSans 224 90 0 0 seg[4]
port 13 nsew signal output
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 seg[5]
port 14 nsew signal output
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 seg[6]
port 15 nsew signal output
rlabel metal1 9982 17408 9982 17408 0 VGND
rlabel metal1 9982 16864 9982 16864 0 VPWR
rlabel metal3 1050 9588 1050 9588 0 net1
rlabel metal3 751 11628 751 11628 0 net10
rlabel metal3 751 8908 751 8908 0 net11
rlabel metal3 1050 10948 1050 10948 0 net2
rlabel metal2 18538 10353 18538 10353 0 net3
rlabel metal2 9706 1588 9706 1588 0 net4
rlabel metal1 9752 17170 9752 17170 0 net5
rlabel metal1 10304 17170 10304 17170 0 net6
rlabel metal3 751 10268 751 10268 0 net7
rlabel metal2 10350 1027 10350 1027 0 net8
rlabel metal3 1050 8228 1050 8228 0 net9
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
