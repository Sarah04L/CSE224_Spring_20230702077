VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO myBasic_ALU
  CLASS BLOCK ;
  FOREIGN myBasic_ALU ;
  ORIGIN 0.000 0.000 ;
  SIZE 68.230 BY 78.950 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 74.950 22.910 78.950 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 74.950 32.570 78.950 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 64.230 27.240 68.230 27.840 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END A[7]
  PIN B[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END B[0]
  PIN B[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END B[1]
  PIN B[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 74.950 35.790 78.950 ;
    END
  END B[2]
  PIN B[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 74.950 39.010 78.950 ;
    END
  END B[3]
  PIN B[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 64.230 34.040 68.230 34.640 ;
    END
  END B[4]
  PIN B[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END B[5]
  PIN B[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END B[6]
  PIN B[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END B[7]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 15.150 10.640 16.750 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.410 10.640 31.010 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.670 10.640 45.270 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.930 10.640 59.530 68.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 20.520 62.800 22.120 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 34.800 62.800 36.400 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 49.080 62.800 50.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 63.360 62.800 64.960 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 11.850 10.640 13.450 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 26.110 10.640 27.710 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.370 10.640 41.970 68.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.630 10.640 56.230 68.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 17.220 62.800 18.820 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 31.500 62.800 33.100 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 45.780 62.800 47.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 60.060 62.800 61.660 ;
    END
  END VPWR
  PIN opcode[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END opcode[0]
  PIN opcode[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END opcode[1]
  PIN opcode[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END opcode[2]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 64.230 44.240 68.230 44.840 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 64.230 30.640 68.230 31.240 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 64.230 23.840 68.230 24.440 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891000 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END out[8]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 62.750 68.190 ;
      LAYER li1 ;
        RECT 5.520 10.795 62.560 68.085 ;
      LAYER met1 ;
        RECT 4.210 10.640 62.560 68.240 ;
      LAYER met2 ;
        RECT 4.230 74.670 22.350 74.950 ;
        RECT 23.190 74.670 32.010 74.950 ;
        RECT 32.850 74.670 35.230 74.950 ;
        RECT 36.070 74.670 38.450 74.950 ;
        RECT 39.290 74.670 61.090 74.950 ;
        RECT 4.230 4.280 61.090 74.670 ;
        RECT 4.230 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 61.090 4.280 ;
      LAYER met3 ;
        RECT 3.990 62.240 64.230 68.165 ;
        RECT 4.400 60.840 64.230 62.240 ;
        RECT 3.990 58.840 64.230 60.840 ;
        RECT 4.400 57.440 64.230 58.840 ;
        RECT 3.990 55.440 64.230 57.440 ;
        RECT 4.400 54.040 64.230 55.440 ;
        RECT 3.990 45.240 64.230 54.040 ;
        RECT 4.400 43.840 63.830 45.240 ;
        RECT 3.990 41.840 64.230 43.840 ;
        RECT 4.400 40.440 64.230 41.840 ;
        RECT 3.990 38.440 64.230 40.440 ;
        RECT 4.400 37.040 64.230 38.440 ;
        RECT 3.990 35.040 64.230 37.040 ;
        RECT 4.400 33.640 63.830 35.040 ;
        RECT 3.990 31.640 64.230 33.640 ;
        RECT 4.400 30.240 63.830 31.640 ;
        RECT 3.990 28.240 64.230 30.240 ;
        RECT 4.400 26.840 63.830 28.240 ;
        RECT 3.990 24.840 64.230 26.840 ;
        RECT 4.400 23.440 63.830 24.840 ;
        RECT 3.990 10.715 64.230 23.440 ;
  END
END myBasic_ALU
END LIBRARY

