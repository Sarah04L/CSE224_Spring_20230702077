magic
tech sky130A
magscale 1 2
timestamp 1749470101
<< nwell >>
rect 1066 2159 18898 17425
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 842 2128 18860 17456
<< metal2 >>
rect 9678 19200 9734 20000
rect 10322 19200 10378 20000
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 9678 0 9734 800
rect 10322 0 10378 800
<< obsm2 >>
rect 846 19144 9622 19200
rect 9790 19144 10266 19200
rect 10434 19144 18566 19200
rect 846 856 18566 19144
rect 846 800 1250 856
rect 1418 800 9622 856
rect 9790 800 10266 856
rect 10434 800 18566 856
<< metal3 >>
rect 0 11568 800 11688
rect 0 10888 800 11008
rect 0 10208 800 10328
rect 19200 10208 20000 10328
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 0 8168 800 8288
<< obsm3 >>
rect 798 11768 19200 17441
rect 880 11488 19200 11768
rect 798 11088 19200 11488
rect 880 10808 19200 11088
rect 798 10408 19200 10808
rect 880 10128 19120 10408
rect 798 9728 19200 10128
rect 880 9448 19200 9728
rect 798 9048 19200 9448
rect 880 8768 19200 9048
rect 798 8368 19200 8768
rect 880 8088 19200 8368
rect 798 2143 19200 8088
<< metal4 >>
rect 1544 2128 1864 17456
rect 2204 2128 2524 17456
rect 5544 2128 5864 17456
rect 6204 2128 6524 17456
rect 9544 2128 9864 17456
rect 10204 2128 10524 17456
rect 13544 2128 13864 17456
rect 14204 2128 14524 17456
rect 17544 2128 17864 17456
rect 18204 2128 18524 17456
<< metal5 >>
rect 1056 15276 18908 15596
rect 1056 14616 18908 14936
rect 1056 11276 18908 11596
rect 1056 10616 18908 10936
rect 1056 7276 18908 7596
rect 1056 6616 18908 6936
rect 1056 3276 18908 3596
rect 1056 2616 18908 2936
<< labels >>
rlabel metal4 s 2204 2128 2524 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6204 2128 6524 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 10204 2128 10524 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 14204 2128 14524 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 18204 2128 18524 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3276 18908 3596 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7276 18908 7596 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 11276 18908 11596 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 15276 18908 15596 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1544 2128 1864 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5544 2128 5864 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 9544 2128 9864 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 13544 2128 13864 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 17544 2128 17864 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2616 18908 2936 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 6616 18908 6936 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 10616 18908 10936 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 14616 18908 14936 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 9528 800 9648 6 an[0]
port 3 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 an[1]
port 4 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 an[2]
port 5 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 an[3]
port 6 nsew signal output
rlabel metal2 s 18 0 74 800 6 clk
port 7 nsew signal input
rlabel metal2 s 662 0 718 800 6 control
port 8 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 reset
port 9 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 seg[0]
port 10 nsew signal output
rlabel metal3 s 19200 10208 20000 10328 6 seg[1]
port 11 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 seg[2]
port 12 nsew signal output
rlabel metal2 s 9678 19200 9734 20000 6 seg[3]
port 13 nsew signal output
rlabel metal2 s 10322 19200 10378 20000 6 seg[4]
port 14 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 seg[5]
port 15 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 seg[6]
port 16 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 243210
string GDS_FILE /openlane/designs/cpu_lab6/runs/RUN_2025.06.09_11.54.21/results/signoff/cpu_lab6.magic.gds
string GDS_START 23748
<< end >>

