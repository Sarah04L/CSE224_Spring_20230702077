magic
tech sky130A
magscale 1 2
timestamp 1746361102
<< viali >>
rect 7849 13345 7883 13379
rect 4629 13277 4663 13311
rect 6561 13277 6595 13311
rect 7205 13277 7239 13311
rect 8125 13277 8159 13311
rect 4813 13141 4847 13175
rect 6745 13141 6779 13175
rect 7389 13141 7423 13175
rect 1409 12801 1443 12835
rect 4721 12801 4755 12835
rect 5457 12801 5491 12835
rect 6837 12801 6871 12835
rect 7849 12801 7883 12835
rect 9045 12801 9079 12835
rect 4813 12733 4847 12767
rect 5089 12733 5123 12767
rect 5365 12733 5399 12767
rect 6745 12733 6779 12767
rect 7941 12733 7975 12767
rect 9137 12733 9171 12767
rect 8217 12665 8251 12699
rect 9413 12665 9447 12699
rect 1593 12597 1627 12631
rect 5733 12597 5767 12631
rect 7113 12597 7147 12631
rect 4721 12393 4755 12427
rect 4997 12393 5031 12427
rect 5365 12393 5399 12427
rect 7113 12393 7147 12427
rect 8125 12393 8159 12427
rect 9045 12393 9079 12427
rect 9413 12393 9447 12427
rect 9689 12393 9723 12427
rect 5825 12325 5859 12359
rect 10701 12325 10735 12359
rect 2513 12257 2547 12291
rect 2789 12257 2823 12291
rect 5181 12257 5215 12291
rect 5549 12257 5583 12291
rect 6009 12257 6043 12291
rect 6469 12257 6503 12291
rect 6561 12257 6595 12291
rect 6745 12257 6779 12291
rect 6929 12257 6963 12291
rect 10241 12257 10275 12291
rect 2421 12189 2455 12223
rect 2881 12189 2915 12223
rect 2973 12189 3007 12223
rect 3400 12189 3434 12223
rect 4629 12189 4663 12223
rect 4813 12189 4847 12223
rect 4905 12189 4939 12223
rect 5273 12189 5307 12223
rect 5457 12189 5491 12223
rect 6653 12189 6687 12223
rect 7021 12189 7055 12223
rect 7205 12189 7239 12223
rect 8033 12189 8067 12223
rect 8953 12189 8987 12223
rect 10333 12189 10367 12223
rect 10793 12189 10827 12223
rect 10977 12189 11011 12223
rect 9505 12121 9539 12155
rect 3341 12053 3375 12087
rect 3525 12053 3559 12087
rect 5181 12053 5215 12087
rect 8493 12053 8527 12087
rect 9705 12053 9739 12087
rect 9873 12053 9907 12087
rect 10977 12053 11011 12087
rect 1593 11849 1627 11883
rect 3065 11849 3099 11883
rect 3893 11849 3927 11883
rect 4721 11849 4755 11883
rect 4813 11849 4847 11883
rect 4997 11849 5031 11883
rect 7665 11849 7699 11883
rect 7941 11849 7975 11883
rect 9321 11849 9355 11883
rect 9137 11781 9171 11815
rect 1409 11713 1443 11747
rect 3249 11713 3283 11747
rect 3341 11713 3375 11747
rect 3801 11713 3835 11747
rect 3985 11713 4019 11747
rect 4629 11713 4663 11747
rect 7297 11713 7331 11747
rect 7481 11713 7515 11747
rect 7757 11713 7791 11747
rect 7941 11713 7975 11747
rect 8309 11713 8343 11747
rect 9413 11713 9447 11747
rect 9689 11713 9723 11747
rect 9965 11713 9999 11747
rect 10149 11713 10183 11747
rect 10241 11713 10275 11747
rect 10425 11713 10459 11747
rect 3709 11645 3743 11679
rect 4997 11645 5031 11679
rect 8401 11645 8435 11679
rect 8677 11645 8711 11679
rect 9137 11577 9171 11611
rect 9505 11509 9539 11543
rect 10425 11509 10459 11543
rect 2789 11305 2823 11339
rect 3065 11305 3099 11339
rect 3801 11305 3835 11339
rect 5181 11305 5215 11339
rect 5733 11305 5767 11339
rect 6469 11305 6503 11339
rect 7113 11305 7147 11339
rect 8493 11305 8527 11339
rect 10885 11305 10919 11339
rect 1593 11237 1627 11271
rect 6653 11237 6687 11271
rect 7297 11237 7331 11271
rect 6745 11169 6779 11203
rect 7573 11169 7607 11203
rect 10701 11169 10735 11203
rect 11345 11169 11379 11203
rect 11529 11169 11563 11203
rect 1409 11101 1443 11135
rect 3249 11101 3283 11135
rect 3433 11101 3467 11135
rect 3985 11101 4019 11135
rect 4353 11101 4387 11135
rect 4629 11101 4663 11135
rect 4997 11101 5031 11135
rect 5329 11101 5363 11135
rect 5457 11101 5491 11135
rect 7665 11101 7699 11135
rect 7757 11101 7791 11135
rect 7849 11101 7883 11135
rect 8033 11101 8067 11135
rect 8401 11101 8435 11135
rect 8585 11101 8619 11135
rect 10609 11101 10643 11135
rect 11069 11101 11103 11135
rect 2605 11033 2639 11067
rect 2821 11033 2855 11067
rect 4077 11033 4111 11067
rect 4169 11033 4203 11067
rect 4813 11033 4847 11067
rect 4905 11033 4939 11067
rect 5549 11033 5583 11067
rect 5733 11033 5767 11067
rect 6285 11033 6319 11067
rect 6490 11033 6524 11067
rect 11161 11033 11195 11067
rect 2973 10965 3007 10999
rect 7113 10965 7147 10999
rect 7389 10965 7423 10999
rect 8217 10965 8251 10999
rect 4353 10761 4387 10795
rect 7389 10761 7423 10795
rect 2513 10693 2547 10727
rect 6653 10693 6687 10727
rect 2421 10625 2455 10659
rect 2697 10625 2731 10659
rect 3525 10625 3559 10659
rect 3801 10625 3835 10659
rect 3985 10625 4019 10659
rect 4537 10625 4571 10659
rect 4905 10625 4939 10659
rect 7205 10625 7239 10659
rect 10333 10625 10367 10659
rect 10517 10625 10551 10659
rect 10977 10625 11011 10659
rect 3341 10557 3375 10591
rect 4721 10557 4755 10591
rect 10149 10557 10183 10591
rect 10885 10557 10919 10591
rect 3709 10489 3743 10523
rect 2881 10421 2915 10455
rect 4169 10421 4203 10455
rect 5089 10421 5123 10455
rect 6745 10421 6779 10455
rect 11345 10421 11379 10455
rect 2973 10217 3007 10251
rect 10885 10217 10919 10251
rect 2605 10149 2639 10183
rect 7113 10149 7147 10183
rect 10977 10149 11011 10183
rect 11069 10081 11103 10115
rect 6837 10013 6871 10047
rect 7113 10013 7147 10047
rect 10241 10013 10275 10047
rect 10517 10013 10551 10047
rect 10701 10013 10735 10047
rect 10793 10013 10827 10047
rect 2973 9945 3007 9979
rect 3157 9877 3191 9911
rect 6929 9877 6963 9911
rect 10425 9877 10459 9911
rect 5457 9673 5491 9707
rect 7021 9673 7055 9707
rect 7205 9673 7239 9707
rect 2237 9605 2271 9639
rect 4813 9605 4847 9639
rect 7389 9605 7423 9639
rect 2148 9559 2182 9593
rect 2421 9537 2455 9571
rect 3157 9537 3191 9571
rect 3249 9537 3283 9571
rect 5365 9537 5399 9571
rect 5641 9537 5675 9571
rect 6193 9537 6227 9571
rect 6837 9537 6871 9571
rect 7573 9537 7607 9571
rect 7665 9537 7699 9571
rect 8033 9537 8067 9571
rect 8125 9537 8159 9571
rect 8309 9537 8343 9571
rect 2605 9469 2639 9503
rect 2973 9469 3007 9503
rect 3065 9469 3099 9503
rect 5273 9469 5307 9503
rect 5917 9469 5951 9503
rect 6929 9469 6963 9503
rect 7297 9469 7331 9503
rect 5089 9401 5123 9435
rect 7481 9401 7515 9435
rect 2789 9333 2823 9367
rect 5825 9333 5859 9367
rect 6009 9333 6043 9367
rect 6101 9333 6135 9367
rect 6653 9333 6687 9367
rect 8309 9333 8343 9367
rect 2053 9129 2087 9163
rect 3249 9129 3283 9163
rect 4261 9129 4295 9163
rect 5549 9129 5583 9163
rect 8493 9129 8527 9163
rect 11069 9129 11103 9163
rect 1869 9061 1903 9095
rect 3893 9061 3927 9095
rect 4997 9061 5031 9095
rect 11161 9061 11195 9095
rect 1501 8993 1535 9027
rect 3341 8993 3375 9027
rect 6837 8993 6871 9027
rect 7113 8993 7147 9027
rect 9229 8993 9263 9027
rect 9505 8993 9539 9027
rect 10517 8993 10551 9027
rect 10701 8993 10735 9027
rect 2237 8925 2271 8959
rect 2329 8925 2363 8959
rect 2513 8925 2547 8959
rect 2605 8925 2639 8959
rect 2822 8925 2856 8959
rect 3433 8925 3467 8959
rect 3617 8925 3651 8959
rect 3801 8925 3835 8959
rect 4077 8925 4111 8959
rect 5178 8925 5212 8959
rect 5641 8925 5675 8959
rect 6745 8925 6779 8959
rect 7849 8925 7883 8959
rect 7941 8925 7975 8959
rect 8217 8925 8251 8959
rect 8309 8925 8343 8959
rect 9137 8925 9171 8959
rect 9781 8925 9815 8959
rect 9873 8925 9907 8959
rect 10425 8925 10459 8959
rect 10793 8925 10827 8959
rect 11069 8925 11103 8959
rect 11437 8925 11471 8959
rect 11897 8925 11931 8959
rect 2947 8857 2981 8891
rect 8125 8857 8159 8891
rect 10333 8857 10367 8891
rect 10885 8857 10919 8891
rect 11161 8857 11195 8891
rect 1961 8789 1995 8823
rect 2697 8789 2731 8823
rect 3433 8789 3467 8823
rect 5181 8789 5215 8823
rect 10701 8789 10735 8823
rect 11345 8789 11379 8823
rect 12081 8789 12115 8823
rect 2145 8585 2179 8619
rect 3985 8585 4019 8619
rect 4169 8585 4203 8619
rect 8033 8585 8067 8619
rect 9873 8585 9907 8619
rect 11345 8585 11379 8619
rect 11529 8585 11563 8619
rect 1685 8517 1719 8551
rect 1901 8517 1935 8551
rect 2697 8517 2731 8551
rect 5181 8517 5215 8551
rect 5273 8517 5307 8551
rect 9689 8517 9723 8551
rect 2329 8449 2363 8483
rect 3157 8449 3191 8483
rect 3433 8449 3467 8483
rect 3801 8449 3835 8483
rect 4353 8449 4387 8483
rect 4445 8449 4479 8483
rect 4721 8449 4755 8483
rect 4905 8449 4939 8483
rect 4997 8449 5031 8483
rect 5365 8449 5399 8483
rect 5825 8449 5859 8483
rect 5917 8449 5951 8483
rect 6193 8449 6227 8483
rect 8217 8449 8251 8483
rect 8309 8449 8343 8483
rect 8585 8449 8619 8483
rect 9321 8449 9355 8483
rect 9505 8449 9539 8483
rect 9781 8449 9815 8483
rect 9965 8449 9999 8483
rect 10885 8449 10919 8483
rect 11069 8449 11103 8483
rect 11161 8449 11195 8483
rect 11805 8449 11839 8483
rect 2605 8381 2639 8415
rect 3341 8381 3375 8415
rect 5641 8381 5675 8415
rect 6101 8381 6135 8415
rect 11529 8381 11563 8415
rect 2053 8313 2087 8347
rect 4629 8313 4663 8347
rect 8493 8313 8527 8347
rect 10977 8313 11011 8347
rect 11713 8313 11747 8347
rect 1869 8245 1903 8279
rect 2513 8245 2547 8279
rect 5549 8245 5583 8279
rect 1869 8041 1903 8075
rect 2605 8041 2639 8075
rect 4813 8041 4847 8075
rect 5457 8041 5491 8075
rect 7941 8041 7975 8075
rect 10885 8041 10919 8075
rect 1501 7973 1535 8007
rect 2789 7973 2823 8007
rect 10977 7973 11011 8007
rect 7481 7905 7515 7939
rect 1685 7837 1719 7871
rect 2053 7837 2087 7871
rect 2329 7837 2363 7871
rect 2605 7837 2639 7871
rect 2697 7837 2731 7871
rect 2881 7837 2915 7871
rect 4537 7837 4571 7871
rect 5181 7837 5215 7871
rect 5273 7837 5307 7871
rect 6745 7837 6779 7871
rect 7573 7837 7607 7871
rect 10333 7837 10367 7871
rect 10425 7837 10459 7871
rect 11805 7837 11839 7871
rect 2421 7769 2455 7803
rect 4629 7769 4663 7803
rect 4813 7769 4847 7803
rect 5457 7769 5491 7803
rect 10609 7769 10643 7803
rect 11345 7769 11379 7803
rect 11621 7769 11655 7803
rect 7205 7701 7239 7735
rect 11437 7701 11471 7735
rect 1961 7497 1995 7531
rect 6561 7497 6595 7531
rect 7757 7497 7791 7531
rect 11713 7497 11747 7531
rect 2329 7429 2363 7463
rect 2881 7429 2915 7463
rect 3065 7429 3099 7463
rect 4997 7429 5031 7463
rect 10333 7429 10367 7463
rect 10517 7429 10551 7463
rect 1685 7361 1719 7395
rect 1777 7361 1811 7395
rect 2513 7361 2547 7395
rect 2789 7361 2823 7395
rect 3341 7361 3375 7395
rect 5181 7361 5215 7395
rect 5457 7361 5491 7395
rect 6377 7361 6411 7395
rect 6561 7361 6595 7395
rect 6929 7361 6963 7395
rect 7389 7361 7423 7395
rect 7941 7361 7975 7395
rect 8217 7361 8251 7395
rect 10701 7361 10735 7395
rect 10977 7361 11011 7395
rect 11161 7361 11195 7395
rect 11529 7361 11563 7395
rect 11805 7361 11839 7395
rect 5365 7293 5399 7327
rect 6653 7293 6687 7327
rect 7113 7293 7147 7327
rect 7297 7293 7331 7327
rect 8125 7293 8159 7327
rect 11253 7293 11287 7327
rect 3249 7225 3283 7259
rect 5641 7225 5675 7259
rect 6745 7225 6779 7259
rect 8033 7225 8067 7259
rect 11529 7225 11563 7259
rect 1501 7157 1535 7191
rect 2697 7157 2731 7191
rect 2789 7157 2823 7191
rect 8401 7157 8435 7191
rect 10793 7157 10827 7191
rect 2145 6953 2179 6987
rect 7481 6953 7515 6987
rect 7573 6885 7607 6919
rect 8401 6817 8435 6851
rect 10609 6817 10643 6851
rect 12173 6817 12207 6851
rect 2329 6749 2363 6783
rect 2697 6749 2731 6783
rect 3065 6749 3099 6783
rect 3157 6749 3191 6783
rect 3249 6749 3283 6783
rect 3433 6749 3467 6783
rect 5181 6749 5215 6783
rect 7389 6749 7423 6783
rect 7665 6749 7699 6783
rect 7849 6749 7883 6783
rect 8309 6749 8343 6783
rect 9781 6749 9815 6783
rect 9965 6749 9999 6783
rect 10057 6749 10091 6783
rect 10701 6749 10735 6783
rect 11069 6749 11103 6783
rect 11253 6749 11287 6783
rect 11897 6749 11931 6783
rect 2421 6681 2455 6715
rect 2513 6681 2547 6715
rect 2789 6613 2823 6647
rect 5365 6613 5399 6647
rect 7113 6613 7147 6647
rect 8677 6613 8711 6647
rect 9597 6613 9631 6647
rect 2605 6409 2639 6443
rect 3525 6409 3559 6443
rect 8677 6409 8711 6443
rect 10977 6409 11011 6443
rect 11345 6409 11379 6443
rect 10793 6341 10827 6375
rect 11989 6341 12023 6375
rect 1501 6273 1535 6307
rect 2789 6273 2823 6307
rect 3065 6273 3099 6307
rect 3433 6273 3467 6307
rect 3525 6273 3559 6307
rect 3801 6273 3835 6307
rect 4077 6273 4111 6307
rect 5089 6273 5123 6307
rect 5181 6273 5215 6307
rect 5447 6273 5481 6307
rect 5549 6273 5583 6307
rect 5733 6273 5767 6307
rect 5825 6273 5859 6307
rect 8033 6273 8067 6307
rect 8125 6273 8159 6307
rect 8309 6273 8343 6307
rect 8401 6273 8435 6307
rect 8493 6273 8527 6307
rect 8953 6273 8987 6307
rect 9045 6273 9079 6307
rect 9321 6273 9355 6307
rect 9597 6273 9631 6307
rect 9781 6273 9815 6307
rect 9873 6273 9907 6307
rect 9965 6273 9999 6307
rect 10517 6273 10551 6307
rect 10609 6273 10643 6307
rect 10885 6273 10919 6307
rect 11161 6273 11195 6307
rect 2881 6205 2915 6239
rect 2973 6205 3007 6239
rect 4905 6205 4939 6239
rect 4997 6205 5031 6239
rect 5365 6205 5399 6239
rect 10425 6205 10459 6239
rect 11529 6205 11563 6239
rect 3801 6137 3835 6171
rect 9229 6137 9263 6171
rect 11621 6137 11655 6171
rect 1777 6069 1811 6103
rect 6009 6069 6043 6103
rect 8769 6069 8803 6103
rect 9781 6069 9815 6103
rect 10793 6069 10827 6103
rect 2421 5865 2455 5899
rect 3157 5865 3191 5899
rect 3341 5865 3375 5899
rect 5641 5865 5675 5899
rect 5825 5865 5859 5899
rect 8493 5865 8527 5899
rect 11069 5865 11103 5899
rect 2789 5797 2823 5831
rect 4997 5797 5031 5831
rect 6285 5797 6319 5831
rect 4353 5729 4387 5763
rect 11897 5729 11931 5763
rect 1685 5661 1719 5695
rect 2053 5661 2087 5695
rect 2605 5661 2639 5695
rect 2789 5661 2823 5695
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 4261 5661 4295 5695
rect 4445 5661 4479 5695
rect 4721 5661 4755 5695
rect 4813 5661 4847 5695
rect 5214 5661 5248 5695
rect 5733 5661 5767 5695
rect 6009 5661 6043 5695
rect 6101 5661 6135 5695
rect 6377 5661 6411 5695
rect 7205 5661 7239 5695
rect 7297 5661 7331 5695
rect 7481 5661 7515 5695
rect 7573 5661 7607 5695
rect 8217 5661 8251 5695
rect 8309 5661 8343 5695
rect 10425 5661 10459 5695
rect 10517 5661 10551 5695
rect 10701 5661 10735 5695
rect 10793 5661 10827 5695
rect 11069 5661 11103 5695
rect 11253 5661 11287 5695
rect 12173 5661 12207 5695
rect 1501 5593 1535 5627
rect 2237 5593 2271 5627
rect 2973 5593 3007 5627
rect 4169 5593 4203 5627
rect 4997 5593 5031 5627
rect 8493 5593 8527 5627
rect 3157 5525 3191 5559
rect 5089 5525 5123 5559
rect 5273 5525 5307 5559
rect 7757 5525 7791 5559
rect 10977 5525 11011 5559
rect 2605 5321 2639 5355
rect 7205 5321 7239 5355
rect 8769 5321 8803 5355
rect 12081 5321 12115 5355
rect 1685 5253 1719 5287
rect 5457 5253 5491 5287
rect 1501 5185 1535 5219
rect 2513 5185 2547 5219
rect 3249 5185 3283 5219
rect 3525 5185 3559 5219
rect 4077 5185 4111 5219
rect 5273 5185 5307 5219
rect 7481 5185 7515 5219
rect 7573 5185 7607 5219
rect 8401 5185 8435 5219
rect 11529 5185 11563 5219
rect 11897 5185 11931 5219
rect 3893 5117 3927 5151
rect 4261 5117 4295 5151
rect 4537 5117 4571 5151
rect 6561 5117 6595 5151
rect 7389 5117 7423 5151
rect 7665 5117 7699 5151
rect 8309 5117 8343 5151
rect 8493 5117 8527 5151
rect 8585 5117 8619 5151
rect 7021 4981 7055 5015
rect 11713 4981 11747 5015
rect 2973 4777 3007 4811
rect 4353 4777 4387 4811
rect 4813 4777 4847 4811
rect 7205 4777 7239 4811
rect 8217 4777 8251 4811
rect 10149 4777 10183 4811
rect 10701 4777 10735 4811
rect 10977 4777 11011 4811
rect 8125 4709 8159 4743
rect 8953 4709 8987 4743
rect 4537 4641 4571 4675
rect 7665 4641 7699 4675
rect 8677 4641 8711 4675
rect 11161 4641 11195 4675
rect 2881 4573 2915 4607
rect 3065 4573 3099 4607
rect 4261 4573 4295 4607
rect 4997 4573 5031 4607
rect 5181 4573 5215 4607
rect 7389 4573 7423 4607
rect 7481 4573 7515 4607
rect 7757 4573 7791 4607
rect 7849 4573 7883 4607
rect 7941 4573 7975 4607
rect 8125 4573 8159 4607
rect 8401 4573 8435 4607
rect 8493 4573 8527 4607
rect 8769 4573 8803 4607
rect 9229 4573 9263 4607
rect 10274 4573 10308 4607
rect 10793 4573 10827 4607
rect 10885 4573 10919 4607
rect 8953 4505 8987 4539
rect 9137 4505 9171 4539
rect 5089 4437 5123 4471
rect 10333 4437 10367 4471
rect 11161 4437 11195 4471
rect 8033 4233 8067 4267
rect 4169 4165 4203 4199
rect 5977 4165 6011 4199
rect 6193 4165 6227 4199
rect 9689 4165 9723 4199
rect 3801 4097 3835 4131
rect 4905 4097 4939 4131
rect 5365 4097 5399 4131
rect 7665 4097 7699 4131
rect 8036 4097 8070 4131
rect 9873 4097 9907 4131
rect 10057 4097 10091 4131
rect 10241 4097 10275 4131
rect 10333 4097 10367 4131
rect 10517 4097 10551 4131
rect 10793 4097 10827 4131
rect 11069 4097 11103 4131
rect 11253 4097 11287 4131
rect 11713 4097 11747 4131
rect 11805 4097 11839 4131
rect 4721 4029 4755 4063
rect 4813 4029 4847 4063
rect 4997 4029 5031 4063
rect 5273 4029 5307 4063
rect 5733 4029 5767 4063
rect 7573 4029 7607 4063
rect 11529 4029 11563 4063
rect 5825 3961 5859 3995
rect 10425 3961 10459 3995
rect 10885 3961 10919 3995
rect 10977 3961 11011 3995
rect 4169 3893 4203 3927
rect 4353 3893 4387 3927
rect 4537 3893 4571 3927
rect 6009 3893 6043 3927
rect 8217 3893 8251 3927
rect 9505 3893 9539 3927
rect 4445 3689 4479 3723
rect 4721 3689 4755 3723
rect 5273 3689 5307 3723
rect 6009 3689 6043 3723
rect 9689 3689 9723 3723
rect 4353 3621 4387 3655
rect 9597 3621 9631 3655
rect 5457 3553 5491 3587
rect 5825 3553 5859 3587
rect 5917 3553 5951 3587
rect 6745 3553 6779 3587
rect 7297 3553 7331 3587
rect 8033 3553 8067 3587
rect 8493 3553 8527 3587
rect 9229 3553 9263 3587
rect 4169 3485 4203 3519
rect 4353 3485 4387 3519
rect 4629 3485 4663 3519
rect 4997 3485 5031 3519
rect 5089 3485 5123 3519
rect 5549 3485 5583 3519
rect 6009 3485 6043 3519
rect 6101 3485 6135 3519
rect 6561 3485 6595 3519
rect 6837 3485 6871 3519
rect 7481 3485 7515 3519
rect 7757 3485 7791 3519
rect 8125 3485 8159 3519
rect 10057 3485 10091 3519
rect 10149 3485 10183 3519
rect 10517 3485 10551 3519
rect 10977 3485 11011 3519
rect 11345 3485 11379 3519
rect 6285 3417 6319 3451
rect 9781 3417 9815 3451
rect 6377 3349 6411 3383
rect 7665 3349 7699 3383
rect 5273 3145 5307 3179
rect 5549 3145 5583 3179
rect 5917 3145 5951 3179
rect 7389 3145 7423 3179
rect 9045 3145 9079 3179
rect 9213 3145 9247 3179
rect 10241 3145 10275 3179
rect 10793 3145 10827 3179
rect 7757 3077 7791 3111
rect 9413 3077 9447 3111
rect 4905 3009 4939 3043
rect 5733 3009 5767 3043
rect 6009 3009 6043 3043
rect 6377 3009 6411 3043
rect 7021 3009 7055 3043
rect 7481 3009 7515 3043
rect 7665 3009 7699 3043
rect 7941 3009 7975 3043
rect 8125 3009 8159 3043
rect 8309 3009 8343 3043
rect 9781 3009 9815 3043
rect 10701 3009 10735 3043
rect 10885 3009 10919 3043
rect 10977 3009 11011 3043
rect 4997 2941 5031 2975
rect 6929 2941 6963 2975
rect 7573 2941 7607 2975
rect 8217 2941 8251 2975
rect 8769 2941 8803 2975
rect 11069 2941 11103 2975
rect 6469 2805 6503 2839
rect 9229 2805 9263 2839
rect 10057 2805 10091 2839
rect 6653 2601 6687 2635
rect 8493 2601 8527 2635
rect 10241 2601 10275 2635
rect 4353 2533 4387 2567
rect 5917 2465 5951 2499
rect 7481 2465 7515 2499
rect 9413 2465 9447 2499
rect 4537 2397 4571 2431
rect 4629 2397 4663 2431
rect 6193 2397 6227 2431
rect 7205 2397 7239 2431
rect 8401 2397 8435 2431
rect 8677 2397 8711 2431
rect 9137 2397 9171 2431
rect 10057 2397 10091 2431
rect 4905 2329 4939 2363
rect 6745 2329 6779 2363
rect 8217 2261 8251 2295
<< metal1 >>
rect 1104 13626 12512 13648
rect 1104 13574 2376 13626
rect 2428 13574 2440 13626
rect 2492 13574 2504 13626
rect 2556 13574 2568 13626
rect 2620 13574 2632 13626
rect 2684 13574 5228 13626
rect 5280 13574 5292 13626
rect 5344 13574 5356 13626
rect 5408 13574 5420 13626
rect 5472 13574 5484 13626
rect 5536 13574 8080 13626
rect 8132 13574 8144 13626
rect 8196 13574 8208 13626
rect 8260 13574 8272 13626
rect 8324 13574 8336 13626
rect 8388 13574 10932 13626
rect 10984 13574 10996 13626
rect 11048 13574 11060 13626
rect 11112 13574 11124 13626
rect 11176 13574 11188 13626
rect 11240 13574 12512 13626
rect 1104 13552 12512 13574
rect 7742 13336 7748 13388
rect 7800 13376 7806 13388
rect 7837 13379 7895 13385
rect 7837 13376 7849 13379
rect 7800 13348 7849 13376
rect 7800 13336 7806 13348
rect 7837 13345 7849 13348
rect 7883 13345 7895 13379
rect 7837 13339 7895 13345
rect 4522 13268 4528 13320
rect 4580 13308 4586 13320
rect 4617 13311 4675 13317
rect 4617 13308 4629 13311
rect 4580 13280 4629 13308
rect 4580 13268 4586 13280
rect 4617 13277 4629 13280
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6512 13280 6561 13308
rect 6512 13268 6518 13280
rect 6549 13277 6561 13280
rect 6595 13277 6607 13311
rect 6549 13271 6607 13277
rect 7098 13268 7104 13320
rect 7156 13308 7162 13320
rect 7193 13311 7251 13317
rect 7193 13308 7205 13311
rect 7156 13280 7205 13308
rect 7156 13268 7162 13280
rect 7193 13277 7205 13280
rect 7239 13277 7251 13311
rect 8113 13311 8171 13317
rect 8113 13308 8125 13311
rect 7193 13271 7251 13277
rect 7852 13280 8125 13308
rect 7852 13252 7880 13280
rect 8113 13277 8125 13280
rect 8159 13277 8171 13311
rect 8113 13271 8171 13277
rect 7834 13200 7840 13252
rect 7892 13200 7898 13252
rect 4614 13132 4620 13184
rect 4672 13172 4678 13184
rect 4801 13175 4859 13181
rect 4801 13172 4813 13175
rect 4672 13144 4813 13172
rect 4672 13132 4678 13144
rect 4801 13141 4813 13144
rect 4847 13141 4859 13175
rect 4801 13135 4859 13141
rect 6270 13132 6276 13184
rect 6328 13172 6334 13184
rect 6733 13175 6791 13181
rect 6733 13172 6745 13175
rect 6328 13144 6745 13172
rect 6328 13132 6334 13144
rect 6733 13141 6745 13144
rect 6779 13141 6791 13175
rect 6733 13135 6791 13141
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7377 13175 7435 13181
rect 7377 13172 7389 13175
rect 7248 13144 7389 13172
rect 7248 13132 7254 13144
rect 7377 13141 7389 13144
rect 7423 13141 7435 13175
rect 7377 13135 7435 13141
rect 1104 13082 12512 13104
rect 1104 13030 3036 13082
rect 3088 13030 3100 13082
rect 3152 13030 3164 13082
rect 3216 13030 3228 13082
rect 3280 13030 3292 13082
rect 3344 13030 5888 13082
rect 5940 13030 5952 13082
rect 6004 13030 6016 13082
rect 6068 13030 6080 13082
rect 6132 13030 6144 13082
rect 6196 13030 8740 13082
rect 8792 13030 8804 13082
rect 8856 13030 8868 13082
rect 8920 13030 8932 13082
rect 8984 13030 8996 13082
rect 9048 13030 11592 13082
rect 11644 13030 11656 13082
rect 11708 13030 11720 13082
rect 11772 13030 11784 13082
rect 11836 13030 11848 13082
rect 11900 13030 12512 13082
rect 1104 13008 12512 13030
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 4706 12792 4712 12844
rect 4764 12792 4770 12844
rect 4982 12792 4988 12844
rect 5040 12832 5046 12844
rect 5445 12835 5503 12841
rect 5445 12832 5457 12835
rect 5040 12804 5457 12832
rect 5040 12792 5046 12804
rect 5445 12801 5457 12804
rect 5491 12801 5503 12835
rect 5445 12795 5503 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 7098 12832 7104 12844
rect 6871 12804 7104 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7098 12792 7104 12804
rect 7156 12792 7162 12844
rect 7650 12792 7656 12844
rect 7708 12832 7714 12844
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 7708 12804 7849 12832
rect 7708 12792 7714 12804
rect 7837 12801 7849 12804
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 9030 12792 9036 12844
rect 9088 12792 9094 12844
rect 4798 12724 4804 12776
rect 4856 12724 4862 12776
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5353 12767 5411 12773
rect 5353 12764 5365 12767
rect 5123 12736 5365 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5353 12733 5365 12736
rect 5399 12764 5411 12767
rect 5810 12764 5816 12776
rect 5399 12736 5816 12764
rect 5399 12733 5411 12736
rect 5353 12727 5411 12733
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 6733 12767 6791 12773
rect 6733 12733 6745 12767
rect 6779 12733 6791 12767
rect 6733 12727 6791 12733
rect 6748 12640 6776 12727
rect 7926 12724 7932 12776
rect 7984 12724 7990 12776
rect 8938 12764 8944 12776
rect 8220 12736 8944 12764
rect 8220 12705 8248 12736
rect 8938 12724 8944 12736
rect 8996 12764 9002 12776
rect 9125 12767 9183 12773
rect 9125 12764 9137 12767
rect 8996 12736 9137 12764
rect 8996 12724 9002 12736
rect 9125 12733 9137 12736
rect 9171 12733 9183 12767
rect 9125 12727 9183 12733
rect 8205 12699 8263 12705
rect 8205 12665 8217 12699
rect 8251 12665 8263 12699
rect 8205 12659 8263 12665
rect 9401 12699 9459 12705
rect 9401 12665 9413 12699
rect 9447 12696 9459 12699
rect 10318 12696 10324 12708
rect 9447 12668 10324 12696
rect 9447 12665 9459 12668
rect 9401 12659 9459 12665
rect 10318 12656 10324 12668
rect 10376 12656 10382 12708
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 1670 12628 1676 12640
rect 1627 12600 1676 12628
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 1670 12588 1676 12600
rect 1728 12588 1734 12640
rect 5721 12631 5779 12637
rect 5721 12597 5733 12631
rect 5767 12628 5779 12631
rect 6730 12628 6736 12640
rect 5767 12600 6736 12628
rect 5767 12597 5779 12600
rect 5721 12591 5779 12597
rect 6730 12588 6736 12600
rect 6788 12588 6794 12640
rect 7101 12631 7159 12637
rect 7101 12597 7113 12631
rect 7147 12628 7159 12631
rect 10226 12628 10232 12640
rect 7147 12600 10232 12628
rect 7147 12597 7159 12600
rect 7101 12591 7159 12597
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 1104 12538 12512 12560
rect 1104 12486 2376 12538
rect 2428 12486 2440 12538
rect 2492 12486 2504 12538
rect 2556 12486 2568 12538
rect 2620 12486 2632 12538
rect 2684 12486 5228 12538
rect 5280 12486 5292 12538
rect 5344 12486 5356 12538
rect 5408 12486 5420 12538
rect 5472 12486 5484 12538
rect 5536 12486 8080 12538
rect 8132 12486 8144 12538
rect 8196 12486 8208 12538
rect 8260 12486 8272 12538
rect 8324 12486 8336 12538
rect 8388 12486 10932 12538
rect 10984 12486 10996 12538
rect 11048 12486 11060 12538
rect 11112 12486 11124 12538
rect 11176 12486 11188 12538
rect 11240 12486 12512 12538
rect 1104 12464 12512 12486
rect 4706 12384 4712 12436
rect 4764 12384 4770 12436
rect 4798 12384 4804 12436
rect 4856 12424 4862 12436
rect 4985 12427 5043 12433
rect 4985 12424 4997 12427
rect 4856 12396 4997 12424
rect 4856 12384 4862 12396
rect 4985 12393 4997 12396
rect 5031 12424 5043 12427
rect 5353 12427 5411 12433
rect 5353 12424 5365 12427
rect 5031 12396 5365 12424
rect 5031 12393 5043 12396
rect 4985 12387 5043 12393
rect 5353 12393 5365 12396
rect 5399 12393 5411 12427
rect 5353 12387 5411 12393
rect 7098 12384 7104 12436
rect 7156 12384 7162 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 8113 12427 8171 12433
rect 8113 12424 8125 12427
rect 7708 12396 8125 12424
rect 7708 12384 7714 12396
rect 8113 12393 8125 12396
rect 8159 12393 8171 12427
rect 8113 12387 8171 12393
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 9030 12424 9036 12436
rect 8720 12396 9036 12424
rect 8720 12384 8726 12396
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 9674 12424 9680 12436
rect 9447 12396 9680 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 2866 12316 2872 12368
rect 2924 12356 2930 12368
rect 2924 12328 4568 12356
rect 2924 12316 2930 12328
rect 2501 12291 2559 12297
rect 2501 12257 2513 12291
rect 2547 12257 2559 12291
rect 2501 12251 2559 12257
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 3602 12288 3608 12300
rect 2823 12260 3608 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2516 12220 2544 12251
rect 3602 12248 3608 12260
rect 3660 12248 3666 12300
rect 4540 12232 4568 12328
rect 4724 12288 4752 12384
rect 5000 12328 5580 12356
rect 5000 12300 5028 12328
rect 4724 12260 4936 12288
rect 2866 12220 2872 12232
rect 2516 12192 2872 12220
rect 2409 12183 2467 12189
rect 2424 12152 2452 12183
rect 2866 12180 2872 12192
rect 2924 12180 2930 12232
rect 3418 12229 3424 12232
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 2961 12183 3019 12189
rect 3388 12223 3424 12229
rect 3388 12189 3400 12223
rect 3388 12183 3424 12189
rect 2976 12152 3004 12183
rect 3418 12180 3424 12183
rect 3476 12180 3482 12232
rect 4522 12180 4528 12232
rect 4580 12220 4586 12232
rect 4617 12223 4675 12229
rect 4617 12220 4629 12223
rect 4580 12192 4629 12220
rect 4580 12180 4586 12192
rect 4617 12189 4629 12192
rect 4663 12189 4675 12223
rect 4798 12220 4804 12232
rect 4617 12183 4675 12189
rect 4724 12192 4804 12220
rect 3878 12152 3884 12164
rect 2424 12124 3884 12152
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 3970 12112 3976 12164
rect 4028 12152 4034 12164
rect 4724 12152 4752 12192
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 4908 12229 4936 12260
rect 4982 12248 4988 12300
rect 5040 12248 5046 12300
rect 5166 12248 5172 12300
rect 5224 12288 5230 12300
rect 5552 12297 5580 12328
rect 5810 12316 5816 12368
rect 5868 12316 5874 12368
rect 6822 12356 6828 12368
rect 6564 12328 6828 12356
rect 6564 12297 6592 12328
rect 6822 12316 6828 12328
rect 6880 12316 6886 12368
rect 10689 12359 10747 12365
rect 10689 12325 10701 12359
rect 10735 12356 10747 12359
rect 10778 12356 10784 12368
rect 10735 12328 10784 12356
rect 10735 12325 10747 12328
rect 10689 12319 10747 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 5537 12291 5595 12297
rect 5224 12260 5304 12288
rect 5224 12248 5230 12260
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12189 4951 12223
rect 4893 12183 4951 12189
rect 5000 12152 5028 12248
rect 5276 12229 5304 12260
rect 5537 12257 5549 12291
rect 5583 12257 5595 12291
rect 5537 12251 5595 12257
rect 5997 12291 6055 12297
rect 5997 12257 6009 12291
rect 6043 12288 6055 12291
rect 6457 12291 6515 12297
rect 6457 12288 6469 12291
rect 6043 12260 6469 12288
rect 6043 12257 6055 12260
rect 5997 12251 6055 12257
rect 6457 12257 6469 12260
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 6549 12291 6607 12297
rect 6549 12257 6561 12291
rect 6595 12257 6607 12291
rect 6549 12251 6607 12257
rect 6730 12248 6736 12300
rect 6788 12248 6794 12300
rect 6917 12291 6975 12297
rect 6917 12257 6929 12291
rect 6963 12288 6975 12291
rect 10229 12291 10287 12297
rect 10229 12288 10241 12291
rect 6963 12260 10241 12288
rect 6963 12257 6975 12260
rect 6917 12251 6975 12257
rect 10229 12257 10241 12260
rect 10275 12288 10287 12291
rect 10275 12260 10824 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 5445 12223 5503 12229
rect 5445 12189 5457 12223
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 7009 12223 7067 12229
rect 7009 12220 7021 12223
rect 6687 12192 7021 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 7009 12189 7021 12192
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12189 7251 12223
rect 7193 12183 7251 12189
rect 4028 12124 4752 12152
rect 4816 12124 5028 12152
rect 4028 12112 4034 12124
rect 2958 12044 2964 12096
rect 3016 12084 3022 12096
rect 3329 12087 3387 12093
rect 3329 12084 3341 12087
rect 3016 12056 3341 12084
rect 3016 12044 3022 12056
rect 3329 12053 3341 12056
rect 3375 12053 3387 12087
rect 3329 12047 3387 12053
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 4816 12084 4844 12124
rect 5074 12112 5080 12164
rect 5132 12152 5138 12164
rect 5460 12152 5488 12183
rect 5132 12124 5488 12152
rect 5132 12112 5138 12124
rect 5534 12112 5540 12164
rect 5592 12152 5598 12164
rect 6656 12152 6684 12183
rect 5592 12124 6684 12152
rect 5592 12112 5598 12124
rect 6822 12112 6828 12164
rect 6880 12152 6886 12164
rect 7208 12152 7236 12183
rect 7926 12180 7932 12232
rect 7984 12220 7990 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7984 12192 8033 12220
rect 7984 12180 7990 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 6880 12124 7236 12152
rect 6880 12112 6886 12124
rect 3559 12056 4844 12084
rect 5169 12087 5227 12093
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 8036 12084 8064 12183
rect 8938 12180 8944 12232
rect 8996 12180 9002 12232
rect 10318 12180 10324 12232
rect 10376 12180 10382 12232
rect 10796 12229 10824 12260
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12189 10839 12223
rect 10781 12183 10839 12189
rect 10965 12223 11023 12229
rect 10965 12189 10977 12223
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 9493 12155 9551 12161
rect 9493 12121 9505 12155
rect 9539 12121 9551 12155
rect 10336 12152 10364 12180
rect 10980 12152 11008 12183
rect 10336 12124 11008 12152
rect 9493 12115 9551 12121
rect 5215 12056 8064 12084
rect 8481 12087 8539 12093
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 9306 12084 9312 12096
rect 8527 12056 9312 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 9306 12044 9312 12056
rect 9364 12084 9370 12096
rect 9508 12084 9536 12115
rect 9364 12056 9536 12084
rect 9364 12044 9370 12056
rect 9582 12044 9588 12096
rect 9640 12084 9646 12096
rect 9693 12087 9751 12093
rect 9693 12084 9705 12087
rect 9640 12056 9705 12084
rect 9640 12044 9646 12056
rect 9693 12053 9705 12056
rect 9739 12053 9751 12087
rect 9693 12047 9751 12053
rect 9861 12087 9919 12093
rect 9861 12053 9873 12087
rect 9907 12084 9919 12087
rect 9950 12084 9956 12096
rect 9907 12056 9956 12084
rect 9907 12053 9919 12056
rect 9861 12047 9919 12053
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10965 12087 11023 12093
rect 10965 12053 10977 12087
rect 11011 12084 11023 12087
rect 11514 12084 11520 12096
rect 11011 12056 11520 12084
rect 11011 12053 11023 12056
rect 10965 12047 11023 12053
rect 11514 12044 11520 12056
rect 11572 12044 11578 12096
rect 1104 11994 12512 12016
rect 1104 11942 3036 11994
rect 3088 11942 3100 11994
rect 3152 11942 3164 11994
rect 3216 11942 3228 11994
rect 3280 11942 3292 11994
rect 3344 11942 5888 11994
rect 5940 11942 5952 11994
rect 6004 11942 6016 11994
rect 6068 11942 6080 11994
rect 6132 11942 6144 11994
rect 6196 11942 8740 11994
rect 8792 11942 8804 11994
rect 8856 11942 8868 11994
rect 8920 11942 8932 11994
rect 8984 11942 8996 11994
rect 9048 11942 11592 11994
rect 11644 11942 11656 11994
rect 11708 11942 11720 11994
rect 11772 11942 11784 11994
rect 11836 11942 11848 11994
rect 11900 11942 12512 11994
rect 1104 11920 12512 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2774 11880 2780 11892
rect 1627 11852 2780 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2774 11840 2780 11852
rect 2832 11840 2838 11892
rect 2866 11840 2872 11892
rect 2924 11880 2930 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 2924 11852 3065 11880
rect 2924 11840 2930 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 3053 11843 3111 11849
rect 3878 11840 3884 11892
rect 3936 11840 3942 11892
rect 4614 11840 4620 11892
rect 4672 11880 4678 11892
rect 4709 11883 4767 11889
rect 4709 11880 4721 11883
rect 4672 11852 4721 11880
rect 4672 11840 4678 11852
rect 4709 11849 4721 11852
rect 4755 11849 4767 11883
rect 4709 11843 4767 11849
rect 4801 11883 4859 11889
rect 4801 11849 4813 11883
rect 4847 11880 4859 11883
rect 4890 11880 4896 11892
rect 4847 11852 4896 11880
rect 4847 11849 4859 11852
rect 4801 11843 4859 11849
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 4985 11883 5043 11889
rect 4985 11849 4997 11883
rect 5031 11880 5043 11883
rect 5166 11880 5172 11892
rect 5031 11852 5172 11880
rect 5031 11849 5043 11852
rect 4985 11843 5043 11849
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 7650 11840 7656 11892
rect 7708 11840 7714 11892
rect 7929 11883 7987 11889
rect 7929 11849 7941 11883
rect 7975 11880 7987 11883
rect 8662 11880 8668 11892
rect 7975 11852 8668 11880
rect 7975 11849 7987 11852
rect 7929 11843 7987 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 9306 11840 9312 11892
rect 9364 11840 9370 11892
rect 9582 11840 9588 11892
rect 9640 11840 9646 11892
rect 5258 11772 5264 11824
rect 5316 11812 5322 11824
rect 9125 11815 9183 11821
rect 9125 11812 9137 11815
rect 5316 11784 7788 11812
rect 5316 11772 5322 11784
rect 1026 11704 1032 11756
rect 1084 11744 1090 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 1084 11716 1409 11744
rect 1084 11704 1090 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 2958 11704 2964 11756
rect 3016 11744 3022 11756
rect 3237 11747 3295 11753
rect 3237 11744 3249 11747
rect 3016 11716 3249 11744
rect 3016 11704 3022 11716
rect 3237 11713 3249 11716
rect 3283 11713 3295 11747
rect 3237 11707 3295 11713
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 3418 11744 3424 11756
rect 3375 11716 3424 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 3418 11704 3424 11716
rect 3476 11704 3482 11756
rect 3789 11747 3847 11753
rect 3789 11713 3801 11747
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 3694 11636 3700 11688
rect 3752 11636 3758 11688
rect 3804 11676 3832 11707
rect 3970 11704 3976 11756
rect 4028 11704 4034 11756
rect 4062 11704 4068 11756
rect 4120 11744 4126 11756
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4120 11716 4629 11744
rect 4120 11704 4126 11716
rect 4617 11713 4629 11716
rect 4663 11713 4675 11747
rect 5534 11744 5540 11756
rect 4617 11707 4675 11713
rect 4724 11716 5540 11744
rect 4724 11676 4752 11716
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 7282 11744 7288 11756
rect 6696 11716 7288 11744
rect 6696 11704 6702 11716
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 7760 11753 7788 11784
rect 8680 11784 9137 11812
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11713 7527 11747
rect 7469 11707 7527 11713
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 3804 11648 4752 11676
rect 4985 11679 5043 11685
rect 2866 11568 2872 11620
rect 2924 11608 2930 11620
rect 3804 11608 3832 11648
rect 4985 11645 4997 11679
rect 5031 11645 5043 11679
rect 4985 11639 5043 11645
rect 2924 11580 3832 11608
rect 5000 11608 5028 11639
rect 5718 11636 5724 11688
rect 5776 11676 5782 11688
rect 7484 11676 7512 11707
rect 7834 11704 7840 11756
rect 7892 11744 7898 11756
rect 7929 11747 7987 11753
rect 7929 11744 7941 11747
rect 7892 11716 7941 11744
rect 7892 11704 7898 11716
rect 7929 11713 7941 11716
rect 7975 11713 7987 11747
rect 7929 11707 7987 11713
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 5776 11648 7512 11676
rect 5776 11636 5782 11648
rect 7558 11636 7564 11688
rect 7616 11676 7622 11688
rect 8312 11676 8340 11707
rect 7616 11648 8340 11676
rect 8389 11679 8447 11685
rect 7616 11636 7622 11648
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 8478 11676 8484 11688
rect 8435 11648 8484 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 8478 11636 8484 11648
rect 8536 11636 8542 11688
rect 8680 11685 8708 11784
rect 9125 11781 9137 11784
rect 9171 11812 9183 11815
rect 9600 11812 9628 11840
rect 11514 11812 11520 11824
rect 9171 11784 9628 11812
rect 10152 11784 11520 11812
rect 9171 11781 9183 11784
rect 9125 11775 9183 11781
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11744 9459 11747
rect 9582 11744 9588 11756
rect 9447 11716 9588 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 9582 11704 9588 11716
rect 9640 11704 9646 11756
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 6270 11608 6276 11620
rect 5000 11580 6276 11608
rect 2924 11568 2930 11580
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 9125 11611 9183 11617
rect 9125 11577 9137 11611
rect 9171 11608 9183 11611
rect 9692 11608 9720 11707
rect 9950 11704 9956 11756
rect 10008 11704 10014 11756
rect 10152 11753 10180 11784
rect 11514 11772 11520 11784
rect 11572 11772 11578 11824
rect 10137 11747 10195 11753
rect 10137 11713 10149 11747
rect 10183 11713 10195 11747
rect 10137 11707 10195 11713
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11713 10471 11747
rect 10413 11707 10471 11713
rect 9968 11676 9996 11704
rect 10244 11676 10272 11707
rect 9968 11648 10272 11676
rect 10428 11608 10456 11707
rect 9171 11580 10456 11608
rect 9171 11577 9183 11580
rect 9125 11571 9183 11577
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 4338 11540 4344 11552
rect 3016 11512 4344 11540
rect 3016 11500 3022 11512
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 5626 11540 5632 11552
rect 4856 11512 5632 11540
rect 4856 11500 4862 11512
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 7282 11500 7288 11552
rect 7340 11540 7346 11552
rect 7742 11540 7748 11552
rect 7340 11512 7748 11540
rect 7340 11500 7346 11512
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 8570 11500 8576 11552
rect 8628 11540 8634 11552
rect 9493 11543 9551 11549
rect 9493 11540 9505 11543
rect 8628 11512 9505 11540
rect 8628 11500 8634 11512
rect 9493 11509 9505 11512
rect 9539 11509 9551 11543
rect 9493 11503 9551 11509
rect 10413 11543 10471 11549
rect 10413 11509 10425 11543
rect 10459 11540 10471 11543
rect 10594 11540 10600 11552
rect 10459 11512 10600 11540
rect 10459 11509 10471 11512
rect 10413 11503 10471 11509
rect 10594 11500 10600 11512
rect 10652 11500 10658 11552
rect 1104 11450 12512 11472
rect 1104 11398 2376 11450
rect 2428 11398 2440 11450
rect 2492 11398 2504 11450
rect 2556 11398 2568 11450
rect 2620 11398 2632 11450
rect 2684 11398 5228 11450
rect 5280 11398 5292 11450
rect 5344 11398 5356 11450
rect 5408 11398 5420 11450
rect 5472 11398 5484 11450
rect 5536 11398 8080 11450
rect 8132 11398 8144 11450
rect 8196 11398 8208 11450
rect 8260 11398 8272 11450
rect 8324 11398 8336 11450
rect 8388 11398 10932 11450
rect 10984 11398 10996 11450
rect 11048 11398 11060 11450
rect 11112 11398 11124 11450
rect 11176 11398 11188 11450
rect 11240 11398 12512 11450
rect 1104 11376 12512 11398
rect 1670 11296 1676 11348
rect 1728 11336 1734 11348
rect 2406 11336 2412 11348
rect 1728 11308 2412 11336
rect 1728 11296 1734 11308
rect 2406 11296 2412 11308
rect 2464 11336 2470 11348
rect 2777 11339 2835 11345
rect 2777 11336 2789 11339
rect 2464 11308 2789 11336
rect 2464 11296 2470 11308
rect 2777 11305 2789 11308
rect 2823 11336 2835 11339
rect 2866 11336 2872 11348
rect 2823 11308 2872 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3053 11339 3111 11345
rect 3053 11305 3065 11339
rect 3099 11336 3111 11339
rect 3418 11336 3424 11348
rect 3099 11308 3424 11336
rect 3099 11305 3111 11308
rect 3053 11299 3111 11305
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11268 1639 11271
rect 2958 11268 2964 11280
rect 1627 11240 2964 11268
rect 1627 11237 1639 11240
rect 1581 11231 1639 11237
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 2590 11024 2596 11076
rect 2648 11024 2654 11076
rect 2774 11024 2780 11076
rect 2832 11073 2838 11076
rect 2832 11067 2867 11073
rect 2855 11064 2867 11067
rect 3068 11064 3096 11299
rect 3418 11296 3424 11308
rect 3476 11296 3482 11348
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3752 11308 3801 11336
rect 3752 11296 3758 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 3970 11296 3976 11348
rect 4028 11336 4034 11348
rect 4522 11336 4528 11348
rect 4028 11308 4528 11336
rect 4028 11296 4034 11308
rect 4522 11296 4528 11308
rect 4580 11296 4586 11348
rect 5074 11296 5080 11348
rect 5132 11336 5138 11348
rect 5169 11339 5227 11345
rect 5169 11336 5181 11339
rect 5132 11308 5181 11336
rect 5132 11296 5138 11308
rect 5169 11305 5181 11308
rect 5215 11305 5227 11339
rect 5169 11299 5227 11305
rect 5718 11296 5724 11348
rect 5776 11296 5782 11348
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 7006 11336 7012 11348
rect 6503 11308 7012 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 7101 11339 7159 11345
rect 7101 11305 7113 11339
rect 7147 11336 7159 11339
rect 7147 11308 7236 11336
rect 7147 11305 7159 11308
rect 7101 11299 7159 11305
rect 4338 11228 4344 11280
rect 4396 11268 4402 11280
rect 4396 11240 6592 11268
rect 4396 11228 4402 11240
rect 3878 11200 3884 11212
rect 3252 11172 3884 11200
rect 3252 11141 3280 11172
rect 3878 11160 3884 11172
rect 3936 11200 3942 11212
rect 4062 11200 4068 11212
rect 3936 11172 4068 11200
rect 3936 11160 3942 11172
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 6564 11200 6592 11240
rect 6638 11228 6644 11280
rect 6696 11228 6702 11280
rect 7208 11212 7236 11308
rect 8478 11296 8484 11348
rect 8536 11296 8542 11348
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 10873 11339 10931 11345
rect 10873 11336 10885 11339
rect 10744 11308 10885 11336
rect 10744 11296 10750 11308
rect 10873 11305 10885 11308
rect 10919 11305 10931 11339
rect 10873 11299 10931 11305
rect 7285 11271 7343 11277
rect 7285 11237 7297 11271
rect 7331 11268 7343 11271
rect 7331 11240 7604 11268
rect 7331 11237 7343 11240
rect 7285 11231 7343 11237
rect 7576 11212 7604 11240
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 4632 11172 5488 11200
rect 3237 11135 3295 11141
rect 3237 11101 3249 11135
rect 3283 11101 3295 11135
rect 3237 11095 3295 11101
rect 3421 11135 3479 11141
rect 3421 11101 3433 11135
rect 3467 11132 3479 11135
rect 3970 11132 3976 11144
rect 3467 11104 3976 11132
rect 3467 11101 3479 11104
rect 3421 11095 3479 11101
rect 3970 11092 3976 11104
rect 4028 11092 4034 11144
rect 4080 11132 4108 11160
rect 4632 11141 4660 11172
rect 4341 11135 4399 11141
rect 4341 11132 4353 11135
rect 4080 11104 4353 11132
rect 4341 11101 4353 11104
rect 4387 11132 4399 11135
rect 4617 11135 4675 11141
rect 4387 11104 4568 11132
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 2855 11036 3096 11064
rect 2855 11033 2867 11036
rect 2832 11027 2867 11033
rect 2832 11024 2838 11027
rect 3142 11024 3148 11076
rect 3200 11064 3206 11076
rect 4062 11064 4068 11076
rect 3200 11036 4068 11064
rect 3200 11024 3206 11036
rect 4062 11024 4068 11036
rect 4120 11024 4126 11076
rect 4154 11024 4160 11076
rect 4212 11024 4218 11076
rect 2958 10956 2964 11008
rect 3016 10956 3022 11008
rect 4540 10996 4568 11104
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 5460 11141 5488 11172
rect 6564 11172 6745 11200
rect 4985 11135 5043 11141
rect 4985 11132 4997 11135
rect 4764 11104 4997 11132
rect 4764 11092 4770 11104
rect 4985 11101 4997 11104
rect 5031 11101 5043 11135
rect 5317 11135 5375 11141
rect 5317 11132 5329 11135
rect 4985 11095 5043 11101
rect 5092 11104 5329 11132
rect 4801 11067 4859 11073
rect 4801 11033 4813 11067
rect 4847 11033 4859 11067
rect 4801 11027 4859 11033
rect 4816 10996 4844 11027
rect 4890 11024 4896 11076
rect 4948 11064 4954 11076
rect 5092 11064 5120 11104
rect 5317 11101 5329 11104
rect 5363 11101 5375 11135
rect 5317 11095 5375 11101
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 5491 11104 6316 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 6288 11076 6316 11104
rect 4948 11036 5120 11064
rect 5537 11067 5595 11073
rect 4948 11024 4954 11036
rect 5537 11033 5549 11067
rect 5583 11033 5595 11067
rect 5537 11027 5595 11033
rect 4540 10968 4844 10996
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 5552 10996 5580 11027
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 5721 11067 5779 11073
rect 5721 11064 5733 11067
rect 5684 11036 5733 11064
rect 5684 11024 5690 11036
rect 5721 11033 5733 11036
rect 5767 11033 5779 11067
rect 5721 11027 5779 11033
rect 6270 11024 6276 11076
rect 6328 11024 6334 11076
rect 6478 11067 6536 11073
rect 6478 11033 6490 11067
rect 6524 11064 6536 11067
rect 6564 11064 6592 11172
rect 6733 11169 6745 11172
rect 6779 11169 6791 11203
rect 6733 11163 6791 11169
rect 7190 11160 7196 11212
rect 7248 11160 7254 11212
rect 7558 11160 7564 11212
rect 7616 11160 7622 11212
rect 10689 11203 10747 11209
rect 10689 11169 10701 11203
rect 10735 11200 10747 11203
rect 11333 11203 11391 11209
rect 11333 11200 11345 11203
rect 10735 11172 11345 11200
rect 10735 11169 10747 11172
rect 10689 11163 10747 11169
rect 11333 11169 11345 11172
rect 11379 11169 11391 11203
rect 11333 11163 11391 11169
rect 11514 11160 11520 11212
rect 11572 11160 11578 11212
rect 7650 11132 7656 11144
rect 6524 11036 6592 11064
rect 6656 11104 7656 11132
rect 6524 11033 6536 11036
rect 6478 11027 6536 11033
rect 6656 10996 6684 11104
rect 7650 11092 7656 11104
rect 7708 11092 7714 11144
rect 7745 11135 7803 11141
rect 7745 11101 7757 11135
rect 7791 11101 7803 11135
rect 7745 11095 7803 11101
rect 6822 11024 6828 11076
rect 6880 11064 6886 11076
rect 7760 11064 7788 11095
rect 7834 11092 7840 11144
rect 7892 11092 7898 11144
rect 7926 11092 7932 11144
rect 7984 11132 7990 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 7984 11104 8033 11132
rect 7984 11092 7990 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 8389 11135 8447 11141
rect 8389 11101 8401 11135
rect 8435 11101 8447 11135
rect 8389 11095 8447 11101
rect 8404 11064 8432 11095
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 8573 11135 8631 11141
rect 8573 11132 8585 11135
rect 8536 11104 8585 11132
rect 8536 11092 8542 11104
rect 8573 11101 8585 11104
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 10778 11092 10784 11144
rect 10836 11132 10842 11144
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 10836 11104 11069 11132
rect 10836 11092 10842 11104
rect 11057 11101 11069 11104
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 6880 11036 8432 11064
rect 6880 11024 6886 11036
rect 5132 10968 6684 10996
rect 5132 10956 5138 10968
rect 6914 10956 6920 11008
rect 6972 10996 6978 11008
rect 7101 10999 7159 11005
rect 7101 10996 7113 10999
rect 6972 10968 7113 10996
rect 6972 10956 6978 10968
rect 7101 10965 7113 10968
rect 7147 10965 7159 10999
rect 7101 10959 7159 10965
rect 7374 10956 7380 11008
rect 7432 10956 7438 11008
rect 8220 11005 8248 11036
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 11149 11067 11207 11073
rect 11149 11064 11161 11067
rect 10928 11036 11161 11064
rect 10928 11024 10934 11036
rect 11149 11033 11161 11036
rect 11195 11033 11207 11067
rect 11149 11027 11207 11033
rect 8205 10999 8263 11005
rect 8205 10965 8217 10999
rect 8251 10965 8263 10999
rect 8205 10959 8263 10965
rect 1104 10906 12512 10928
rect 1104 10854 3036 10906
rect 3088 10854 3100 10906
rect 3152 10854 3164 10906
rect 3216 10854 3228 10906
rect 3280 10854 3292 10906
rect 3344 10854 5888 10906
rect 5940 10854 5952 10906
rect 6004 10854 6016 10906
rect 6068 10854 6080 10906
rect 6132 10854 6144 10906
rect 6196 10854 8740 10906
rect 8792 10854 8804 10906
rect 8856 10854 8868 10906
rect 8920 10854 8932 10906
rect 8984 10854 8996 10906
rect 9048 10854 11592 10906
rect 11644 10854 11656 10906
rect 11708 10854 11720 10906
rect 11772 10854 11784 10906
rect 11836 10854 11848 10906
rect 11900 10854 12512 10906
rect 1104 10832 12512 10854
rect 4338 10752 4344 10804
rect 4396 10752 4402 10804
rect 4890 10752 4896 10804
rect 4948 10752 4954 10804
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 7190 10792 7196 10804
rect 5684 10764 7196 10792
rect 5684 10752 5690 10764
rect 7190 10752 7196 10764
rect 7248 10792 7254 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 7248 10764 7389 10792
rect 7248 10752 7254 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 7377 10755 7435 10761
rect 1670 10684 1676 10736
rect 1728 10724 1734 10736
rect 2501 10727 2559 10733
rect 2501 10724 2513 10727
rect 1728 10696 2513 10724
rect 1728 10684 1734 10696
rect 2501 10693 2513 10696
rect 2547 10724 2559 10727
rect 2590 10724 2596 10736
rect 2547 10696 2596 10724
rect 2547 10693 2559 10696
rect 2501 10687 2559 10693
rect 2590 10684 2596 10696
rect 2648 10724 2654 10736
rect 4908 10724 4936 10752
rect 2648 10696 4936 10724
rect 2648 10684 2654 10696
rect 6270 10684 6276 10736
rect 6328 10724 6334 10736
rect 6641 10727 6699 10733
rect 6641 10724 6653 10727
rect 6328 10696 6653 10724
rect 6328 10684 6334 10696
rect 6641 10693 6653 10696
rect 6687 10693 6699 10727
rect 6641 10687 6699 10693
rect 10870 10684 10876 10736
rect 10928 10684 10934 10736
rect 1946 10616 1952 10668
rect 2004 10656 2010 10668
rect 2406 10656 2412 10668
rect 2004 10628 2412 10656
rect 2004 10616 2010 10628
rect 2406 10616 2412 10628
rect 2464 10616 2470 10668
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2774 10656 2780 10668
rect 2731 10628 2780 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 2958 10616 2964 10668
rect 3016 10656 3022 10668
rect 3513 10659 3571 10665
rect 3513 10656 3525 10659
rect 3016 10628 3525 10656
rect 3016 10616 3022 10628
rect 3513 10625 3525 10628
rect 3559 10656 3571 10659
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3559 10628 3801 10656
rect 3559 10625 3571 10628
rect 3513 10619 3571 10625
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10588 3387 10591
rect 3602 10588 3608 10600
rect 3375 10560 3608 10588
rect 3375 10557 3387 10560
rect 3329 10551 3387 10557
rect 3602 10548 3608 10560
rect 3660 10588 3666 10600
rect 3988 10588 4016 10619
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4525 10659 4583 10665
rect 4525 10656 4537 10659
rect 4212 10628 4537 10656
rect 4212 10616 4218 10628
rect 4525 10625 4537 10628
rect 4571 10656 4583 10659
rect 4614 10656 4620 10668
rect 4571 10628 4620 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 4614 10616 4620 10628
rect 4672 10656 4678 10668
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4672 10628 4905 10656
rect 4672 10616 4678 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 7064 10628 7205 10656
rect 7064 10616 7070 10628
rect 7193 10625 7205 10628
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 10226 10616 10232 10668
rect 10284 10656 10290 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 10284 10628 10333 10656
rect 10284 10616 10290 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10505 10659 10563 10665
rect 10505 10625 10517 10659
rect 10551 10656 10563 10659
rect 10686 10656 10692 10668
rect 10551 10628 10692 10656
rect 10551 10625 10563 10628
rect 10505 10619 10563 10625
rect 10686 10616 10692 10628
rect 10744 10656 10750 10668
rect 10888 10656 10916 10684
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10744 10628 10977 10656
rect 10744 10616 10750 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 3660 10560 4016 10588
rect 3660 10548 3666 10560
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 4709 10591 4767 10597
rect 4709 10588 4721 10591
rect 4120 10560 4721 10588
rect 4120 10548 4126 10560
rect 4709 10557 4721 10560
rect 4755 10557 4767 10591
rect 4709 10551 4767 10557
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10557 10195 10591
rect 10137 10551 10195 10557
rect 3697 10523 3755 10529
rect 3697 10489 3709 10523
rect 3743 10520 3755 10523
rect 4798 10520 4804 10532
rect 3743 10492 4804 10520
rect 3743 10489 3755 10492
rect 3697 10483 3755 10489
rect 4798 10480 4804 10492
rect 4856 10520 4862 10532
rect 10152 10520 10180 10551
rect 10778 10548 10784 10600
rect 10836 10588 10842 10600
rect 10873 10591 10931 10597
rect 10873 10588 10885 10591
rect 10836 10560 10885 10588
rect 10836 10548 10842 10560
rect 10873 10557 10885 10560
rect 10919 10557 10931 10591
rect 10873 10551 10931 10557
rect 4856 10492 10180 10520
rect 4856 10480 4862 10492
rect 2869 10455 2927 10461
rect 2869 10421 2881 10455
rect 2915 10452 2927 10455
rect 2958 10452 2964 10464
rect 2915 10424 2964 10452
rect 2915 10421 2927 10424
rect 2869 10415 2927 10421
rect 2958 10412 2964 10424
rect 3016 10412 3022 10464
rect 4154 10412 4160 10464
rect 4212 10412 4218 10464
rect 5074 10412 5080 10464
rect 5132 10412 5138 10464
rect 6733 10455 6791 10461
rect 6733 10421 6745 10455
rect 6779 10452 6791 10455
rect 6914 10452 6920 10464
rect 6779 10424 6920 10452
rect 6779 10421 6791 10424
rect 6733 10415 6791 10421
rect 6914 10412 6920 10424
rect 6972 10412 6978 10464
rect 10152 10452 10180 10492
rect 10778 10452 10784 10464
rect 10152 10424 10784 10452
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 11333 10455 11391 10461
rect 11333 10421 11345 10455
rect 11379 10452 11391 10455
rect 11974 10452 11980 10464
rect 11379 10424 11980 10452
rect 11379 10421 11391 10424
rect 11333 10415 11391 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 1104 10362 12512 10384
rect 1104 10310 2376 10362
rect 2428 10310 2440 10362
rect 2492 10310 2504 10362
rect 2556 10310 2568 10362
rect 2620 10310 2632 10362
rect 2684 10310 5228 10362
rect 5280 10310 5292 10362
rect 5344 10310 5356 10362
rect 5408 10310 5420 10362
rect 5472 10310 5484 10362
rect 5536 10310 8080 10362
rect 8132 10310 8144 10362
rect 8196 10310 8208 10362
rect 8260 10310 8272 10362
rect 8324 10310 8336 10362
rect 8388 10310 10932 10362
rect 10984 10310 10996 10362
rect 11048 10310 11060 10362
rect 11112 10310 11124 10362
rect 11176 10310 11188 10362
rect 11240 10310 12512 10362
rect 1104 10288 12512 10310
rect 2961 10251 3019 10257
rect 2961 10217 2973 10251
rect 3007 10248 3019 10251
rect 4706 10248 4712 10260
rect 3007 10220 4712 10248
rect 3007 10217 3019 10220
rect 2961 10211 3019 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 10284 10220 10885 10248
rect 10284 10208 10290 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 2593 10183 2651 10189
rect 2593 10149 2605 10183
rect 2639 10180 2651 10183
rect 2866 10180 2872 10192
rect 2639 10152 2872 10180
rect 2639 10149 2651 10152
rect 2593 10143 2651 10149
rect 2866 10140 2872 10152
rect 2924 10140 2930 10192
rect 7098 10140 7104 10192
rect 7156 10140 7162 10192
rect 10965 10183 11023 10189
rect 10965 10149 10977 10183
rect 11011 10149 11023 10183
rect 10965 10143 11023 10149
rect 10980 10112 11008 10143
rect 10520 10084 11008 10112
rect 11057 10115 11115 10121
rect 6822 10004 6828 10056
rect 6880 10004 6886 10056
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10044 7159 10047
rect 7374 10044 7380 10056
rect 7147 10016 7380 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 7374 10004 7380 10016
rect 7432 10004 7438 10056
rect 10226 10004 10232 10056
rect 10284 10004 10290 10056
rect 10520 10053 10548 10084
rect 11057 10081 11069 10115
rect 11103 10112 11115 10115
rect 11422 10112 11428 10124
rect 11103 10084 11428 10112
rect 11103 10081 11115 10084
rect 11057 10075 11115 10081
rect 11422 10072 11428 10084
rect 11480 10072 11486 10124
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 10778 10004 10784 10056
rect 10836 10004 10842 10056
rect 2958 9936 2964 9988
rect 3016 9936 3022 9988
rect 3145 9911 3203 9917
rect 3145 9877 3157 9911
rect 3191 9908 3203 9911
rect 3418 9908 3424 9920
rect 3191 9880 3424 9908
rect 3191 9877 3203 9880
rect 3145 9871 3203 9877
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7650 9908 7656 9920
rect 6972 9880 7656 9908
rect 6972 9868 6978 9880
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 10413 9911 10471 9917
rect 10413 9877 10425 9911
rect 10459 9908 10471 9911
rect 11330 9908 11336 9920
rect 10459 9880 11336 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 11330 9868 11336 9880
rect 11388 9868 11394 9920
rect 1104 9818 12512 9840
rect 1104 9766 3036 9818
rect 3088 9766 3100 9818
rect 3152 9766 3164 9818
rect 3216 9766 3228 9818
rect 3280 9766 3292 9818
rect 3344 9766 5888 9818
rect 5940 9766 5952 9818
rect 6004 9766 6016 9818
rect 6068 9766 6080 9818
rect 6132 9766 6144 9818
rect 6196 9766 8740 9818
rect 8792 9766 8804 9818
rect 8856 9766 8868 9818
rect 8920 9766 8932 9818
rect 8984 9766 8996 9818
rect 9048 9766 11592 9818
rect 11644 9766 11656 9818
rect 11708 9766 11720 9818
rect 11772 9766 11784 9818
rect 11836 9766 11848 9818
rect 11900 9766 12512 9818
rect 1104 9744 12512 9766
rect 4154 9664 4160 9716
rect 4212 9704 4218 9716
rect 5445 9707 5503 9713
rect 5445 9704 5457 9707
rect 4212 9676 5457 9704
rect 4212 9664 4218 9676
rect 5445 9673 5457 9676
rect 5491 9673 5503 9707
rect 5445 9667 5503 9673
rect 6822 9664 6828 9716
rect 6880 9704 6886 9716
rect 7009 9707 7067 9713
rect 7009 9704 7021 9707
rect 6880 9676 7021 9704
rect 6880 9664 6886 9676
rect 7009 9673 7021 9676
rect 7055 9673 7067 9707
rect 7009 9667 7067 9673
rect 2225 9639 2283 9645
rect 2225 9605 2237 9639
rect 2271 9636 2283 9639
rect 2866 9636 2872 9648
rect 2271 9608 2872 9636
rect 2271 9605 2283 9608
rect 2225 9599 2283 9605
rect 2136 9593 2194 9599
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 4798 9596 4804 9648
rect 4856 9596 4862 9648
rect 7024 9636 7052 9667
rect 7190 9664 7196 9716
rect 7248 9664 7254 9716
rect 7024 9608 7328 9636
rect 2136 9580 2148 9593
rect 2182 9580 2194 9593
rect 2130 9528 2136 9580
rect 2188 9528 2194 9580
rect 2409 9571 2467 9577
rect 2409 9568 2421 9571
rect 2240 9540 2421 9568
rect 2240 9512 2268 9540
rect 2409 9537 2421 9540
rect 2455 9537 2467 9571
rect 2409 9531 2467 9537
rect 3142 9528 3148 9580
rect 3200 9528 3206 9580
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3418 9568 3424 9580
rect 3283 9540 3424 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9568 5687 9571
rect 5718 9568 5724 9580
rect 5675 9540 5724 9568
rect 5675 9537 5687 9540
rect 5629 9531 5687 9537
rect 2222 9460 2228 9512
rect 2280 9460 2286 9512
rect 2590 9460 2596 9512
rect 2648 9460 2654 9512
rect 2961 9503 3019 9509
rect 2961 9500 2973 9503
rect 2884 9472 2973 9500
rect 2884 9432 2912 9472
rect 2961 9469 2973 9472
rect 3007 9469 3019 9503
rect 2961 9463 3019 9469
rect 3050 9460 3056 9512
rect 3108 9460 3114 9512
rect 3160 9500 3188 9528
rect 3970 9500 3976 9512
rect 3160 9472 3976 9500
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 5261 9503 5319 9509
rect 5261 9469 5273 9503
rect 5307 9500 5319 9503
rect 5368 9500 5396 9531
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9568 6239 9571
rect 6825 9571 6883 9577
rect 6825 9568 6837 9571
rect 6227 9540 6837 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 6825 9537 6837 9540
rect 6871 9568 6883 9571
rect 7098 9568 7104 9580
rect 6871 9540 7104 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7300 9568 7328 9608
rect 7374 9596 7380 9648
rect 7432 9596 7438 9648
rect 7742 9636 7748 9648
rect 7576 9608 7748 9636
rect 7576 9577 7604 9608
rect 7742 9596 7748 9608
rect 7800 9636 7806 9648
rect 7800 9608 8064 9636
rect 7800 9596 7806 9608
rect 7561 9571 7619 9577
rect 7561 9568 7573 9571
rect 7300 9540 7573 9568
rect 7561 9537 7573 9540
rect 7607 9537 7619 9571
rect 7561 9531 7619 9537
rect 7650 9528 7656 9580
rect 7708 9528 7714 9580
rect 8036 9577 8064 9608
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9537 8079 9571
rect 8021 9531 8079 9537
rect 8113 9571 8171 9577
rect 8113 9537 8125 9571
rect 8159 9537 8171 9571
rect 8113 9531 8171 9537
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8662 9568 8668 9580
rect 8343 9540 8668 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 5307 9472 5396 9500
rect 5905 9503 5963 9509
rect 5307 9469 5319 9472
rect 5261 9463 5319 9469
rect 5905 9469 5917 9503
rect 5951 9469 5963 9503
rect 5905 9463 5963 9469
rect 3694 9432 3700 9444
rect 2884 9404 3700 9432
rect 3694 9392 3700 9404
rect 3752 9392 3758 9444
rect 4798 9392 4804 9444
rect 4856 9432 4862 9444
rect 5077 9435 5135 9441
rect 5077 9432 5089 9435
rect 4856 9404 5089 9432
rect 4856 9392 4862 9404
rect 5077 9401 5089 9404
rect 5123 9401 5135 9435
rect 5920 9432 5948 9463
rect 6914 9460 6920 9512
rect 6972 9460 6978 9512
rect 7285 9503 7343 9509
rect 7285 9469 7297 9503
rect 7331 9500 7343 9503
rect 7668 9500 7696 9528
rect 8128 9500 8156 9531
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 7331 9472 7604 9500
rect 7668 9472 8156 9500
rect 7331 9469 7343 9472
rect 7285 9463 7343 9469
rect 7469 9435 7527 9441
rect 7469 9432 7481 9435
rect 5920 9404 7481 9432
rect 5077 9395 5135 9401
rect 7469 9401 7481 9404
rect 7515 9401 7527 9435
rect 7469 9395 7527 9401
rect 7576 9432 7604 9472
rect 9122 9432 9128 9444
rect 7576 9404 9128 9432
rect 2774 9324 2780 9376
rect 2832 9324 2838 9376
rect 5810 9324 5816 9376
rect 5868 9324 5874 9376
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 5960 9336 6009 9364
rect 5960 9324 5966 9336
rect 5997 9333 6009 9336
rect 6043 9333 6055 9367
rect 5997 9327 6055 9333
rect 6086 9324 6092 9376
rect 6144 9324 6150 9376
rect 6641 9367 6699 9373
rect 6641 9333 6653 9367
rect 6687 9364 6699 9367
rect 6730 9364 6736 9376
rect 6687 9336 6736 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 6730 9324 6736 9336
rect 6788 9324 6794 9376
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 7576 9364 7604 9404
rect 9122 9392 9128 9404
rect 9180 9392 9186 9444
rect 6880 9336 7604 9364
rect 8297 9367 8355 9373
rect 6880 9324 6886 9336
rect 8297 9333 8309 9367
rect 8343 9364 8355 9367
rect 8478 9364 8484 9376
rect 8343 9336 8484 9364
rect 8343 9333 8355 9336
rect 8297 9327 8355 9333
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 1104 9274 12512 9296
rect 1104 9222 2376 9274
rect 2428 9222 2440 9274
rect 2492 9222 2504 9274
rect 2556 9222 2568 9274
rect 2620 9222 2632 9274
rect 2684 9222 5228 9274
rect 5280 9222 5292 9274
rect 5344 9222 5356 9274
rect 5408 9222 5420 9274
rect 5472 9222 5484 9274
rect 5536 9222 8080 9274
rect 8132 9222 8144 9274
rect 8196 9222 8208 9274
rect 8260 9222 8272 9274
rect 8324 9222 8336 9274
rect 8388 9222 10932 9274
rect 10984 9222 10996 9274
rect 11048 9222 11060 9274
rect 11112 9222 11124 9274
rect 11176 9222 11188 9274
rect 11240 9222 12512 9274
rect 1104 9200 12512 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 3237 9163 3295 9169
rect 3237 9160 3249 9163
rect 2087 9132 3249 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 3237 9129 3249 9132
rect 3283 9129 3295 9163
rect 3237 9123 3295 9129
rect 3344 9132 4016 9160
rect 1857 9095 1915 9101
rect 1857 9061 1869 9095
rect 1903 9092 1915 9095
rect 2130 9092 2136 9104
rect 1903 9064 2136 9092
rect 1903 9061 1915 9064
rect 1857 9055 1915 9061
rect 2130 9052 2136 9064
rect 2188 9092 2194 9104
rect 2406 9092 2412 9104
rect 2188 9064 2412 9092
rect 2188 9052 2194 9064
rect 2406 9052 2412 9064
rect 2464 9052 2470 9104
rect 2774 9092 2780 9104
rect 2700 9064 2780 9092
rect 1486 8984 1492 9036
rect 1544 8984 1550 9036
rect 2700 9024 2728 9064
rect 2774 9052 2780 9064
rect 2832 9052 2838 9104
rect 3344 9092 3372 9132
rect 3252 9064 3372 9092
rect 2958 9024 2964 9036
rect 2516 8996 2728 9024
rect 2825 8996 2964 9024
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2516 8965 2544 8996
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 2188 8928 2237 8956
rect 2188 8916 2194 8928
rect 2225 8925 2237 8928
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8925 2559 8959
rect 2501 8919 2559 8925
rect 2332 8888 2360 8919
rect 2590 8916 2596 8968
rect 2648 8916 2654 8968
rect 2825 8965 2853 8996
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 2810 8959 2868 8965
rect 2810 8925 2822 8959
rect 2856 8925 2868 8959
rect 2810 8919 2868 8925
rect 2935 8891 2993 8897
rect 2332 8860 2820 8888
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8820 2007 8823
rect 2222 8820 2228 8832
rect 1995 8792 2228 8820
rect 1995 8789 2007 8792
rect 1949 8783 2007 8789
rect 2222 8780 2228 8792
rect 2280 8780 2286 8832
rect 2314 8780 2320 8832
rect 2372 8820 2378 8832
rect 2685 8823 2743 8829
rect 2685 8820 2697 8823
rect 2372 8792 2697 8820
rect 2372 8780 2378 8792
rect 2685 8789 2697 8792
rect 2731 8789 2743 8823
rect 2792 8820 2820 8860
rect 2935 8857 2947 8891
rect 2981 8888 2993 8891
rect 3252 8888 3280 9064
rect 3510 9052 3516 9104
rect 3568 9092 3574 9104
rect 3881 9095 3939 9101
rect 3881 9092 3893 9095
rect 3568 9064 3893 9092
rect 3568 9052 3574 9064
rect 3881 9061 3893 9064
rect 3927 9061 3939 9095
rect 3988 9092 4016 9132
rect 4246 9120 4252 9172
rect 4304 9120 4310 9172
rect 5537 9163 5595 9169
rect 5537 9129 5549 9163
rect 5583 9160 5595 9163
rect 5810 9160 5816 9172
rect 5583 9132 5816 9160
rect 5583 9129 5595 9132
rect 5537 9123 5595 9129
rect 5810 9120 5816 9132
rect 5868 9120 5874 9172
rect 8481 9163 8539 9169
rect 8481 9129 8493 9163
rect 8527 9160 8539 9163
rect 10226 9160 10232 9172
rect 8527 9132 10232 9160
rect 8527 9129 8539 9132
rect 8481 9123 8539 9129
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 11057 9163 11115 9169
rect 11057 9129 11069 9163
rect 11103 9160 11115 9163
rect 11103 9132 11928 9160
rect 11103 9129 11115 9132
rect 11057 9123 11115 9129
rect 3988 9064 4292 9092
rect 3881 9055 3939 9061
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 9024 3387 9027
rect 4154 9024 4160 9036
rect 3375 8996 4160 9024
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 4154 8984 4160 8996
rect 4212 8984 4218 9036
rect 4264 9024 4292 9064
rect 4982 9052 4988 9104
rect 5040 9052 5046 9104
rect 6086 9052 6092 9104
rect 6144 9092 6150 9104
rect 8570 9092 8576 9104
rect 6144 9064 8576 9092
rect 6144 9052 6150 9064
rect 6270 9024 6276 9036
rect 4264 8996 6276 9024
rect 3418 8916 3424 8968
rect 3476 8916 3482 8968
rect 3602 8916 3608 8968
rect 3660 8916 3666 8968
rect 3786 8916 3792 8968
rect 3844 8916 3850 8968
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8956 4123 8959
rect 4522 8956 4528 8968
rect 4111 8928 4528 8956
rect 4111 8925 4123 8928
rect 4065 8919 4123 8925
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 5166 8959 5224 8965
rect 5166 8925 5178 8959
rect 5212 8956 5224 8959
rect 5258 8956 5264 8968
rect 5212 8928 5264 8956
rect 5212 8925 5224 8928
rect 5166 8919 5224 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 2981 8860 3280 8888
rect 2981 8857 2993 8860
rect 2935 8851 2993 8857
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 2792 8792 3433 8820
rect 2685 8783 2743 8789
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 5169 8823 5227 8829
rect 5169 8789 5181 8823
rect 5215 8820 5227 8823
rect 5460 8820 5488 8996
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 6840 9033 6868 9064
rect 8570 9052 8576 9064
rect 8628 9052 8634 9104
rect 10318 9052 10324 9104
rect 10376 9092 10382 9104
rect 11149 9095 11207 9101
rect 10376 9064 10824 9092
rect 10376 9052 10382 9064
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 7101 9027 7159 9033
rect 7101 8993 7113 9027
rect 7147 9024 7159 9027
rect 7558 9024 7564 9036
rect 7147 8996 7564 9024
rect 7147 8993 7159 8996
rect 7101 8987 7159 8993
rect 7558 8984 7564 8996
rect 7616 8984 7622 9036
rect 7742 8984 7748 9036
rect 7800 9024 7806 9036
rect 9217 9027 9275 9033
rect 7800 8996 8248 9024
rect 7800 8984 7806 8996
rect 5629 8959 5687 8965
rect 5629 8925 5641 8959
rect 5675 8925 5687 8959
rect 5629 8919 5687 8925
rect 5215 8792 5488 8820
rect 5644 8820 5672 8919
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 7374 8916 7380 8968
rect 7432 8956 7438 8968
rect 7837 8959 7895 8965
rect 7837 8956 7849 8959
rect 7432 8928 7849 8956
rect 7432 8916 7438 8928
rect 7837 8925 7849 8928
rect 7883 8925 7895 8959
rect 7837 8919 7895 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8018 8956 8024 8968
rect 7975 8928 8024 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 8220 8965 8248 8996
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 9398 9024 9404 9036
rect 9263 8996 9404 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 9493 9027 9551 9033
rect 9493 8993 9505 9027
rect 9539 9024 9551 9027
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 9539 8996 10517 9024
rect 9539 8993 9551 8996
rect 9493 8987 9551 8993
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8294 8916 8300 8968
rect 8352 8916 8358 8968
rect 9122 8916 9128 8968
rect 9180 8916 9186 8968
rect 9766 8916 9772 8968
rect 9824 8916 9830 8968
rect 9876 8965 9904 8996
rect 10505 8993 10517 8996
rect 10551 8993 10563 9027
rect 10505 8987 10563 8993
rect 10686 8984 10692 9036
rect 10744 8984 10750 9036
rect 10796 8965 10824 9064
rect 11149 9061 11161 9095
rect 11195 9061 11207 9095
rect 11149 9055 11207 9061
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 9861 8919 9919 8925
rect 9968 8928 10425 8956
rect 7650 8848 7656 8900
rect 7708 8888 7714 8900
rect 8110 8888 8116 8900
rect 7708 8860 8116 8888
rect 7708 8848 7714 8860
rect 8110 8848 8116 8860
rect 8168 8848 8174 8900
rect 9784 8888 9812 8916
rect 9968 8888 9996 8928
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 11057 8959 11115 8965
rect 11057 8925 11069 8959
rect 11103 8956 11115 8959
rect 11164 8956 11192 9055
rect 11103 8928 11192 8956
rect 11103 8925 11115 8928
rect 11057 8919 11115 8925
rect 11330 8916 11336 8968
rect 11388 8956 11394 8968
rect 11900 8965 11928 9132
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11388 8928 11437 8956
rect 11388 8916 11394 8928
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8925 11943 8959
rect 11885 8919 11943 8925
rect 9784 8860 9996 8888
rect 10318 8848 10324 8900
rect 10376 8848 10382 8900
rect 10502 8848 10508 8900
rect 10560 8888 10566 8900
rect 10873 8891 10931 8897
rect 10873 8888 10885 8891
rect 10560 8860 10885 8888
rect 10560 8848 10566 8860
rect 10873 8857 10885 8860
rect 10919 8857 10931 8891
rect 10873 8851 10931 8857
rect 11149 8891 11207 8897
rect 11149 8857 11161 8891
rect 11195 8888 11207 8891
rect 11238 8888 11244 8900
rect 11195 8860 11244 8888
rect 11195 8857 11207 8860
rect 11149 8851 11207 8857
rect 11238 8848 11244 8860
rect 11296 8848 11302 8900
rect 9582 8820 9588 8832
rect 5644 8792 9588 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10689 8823 10747 8829
rect 10689 8820 10701 8823
rect 9824 8792 10701 8820
rect 9824 8780 9830 8792
rect 10689 8789 10701 8792
rect 10735 8789 10747 8823
rect 10689 8783 10747 8789
rect 11333 8823 11391 8829
rect 11333 8789 11345 8823
rect 11379 8820 11391 8823
rect 11514 8820 11520 8832
rect 11379 8792 11520 8820
rect 11379 8789 11391 8792
rect 11333 8783 11391 8789
rect 11514 8780 11520 8792
rect 11572 8780 11578 8832
rect 12066 8780 12072 8832
rect 12124 8780 12130 8832
rect 1104 8730 12512 8752
rect 1104 8678 3036 8730
rect 3088 8678 3100 8730
rect 3152 8678 3164 8730
rect 3216 8678 3228 8730
rect 3280 8678 3292 8730
rect 3344 8678 5888 8730
rect 5940 8678 5952 8730
rect 6004 8678 6016 8730
rect 6068 8678 6080 8730
rect 6132 8678 6144 8730
rect 6196 8678 8740 8730
rect 8792 8678 8804 8730
rect 8856 8678 8868 8730
rect 8920 8678 8932 8730
rect 8984 8678 8996 8730
rect 9048 8678 11592 8730
rect 11644 8678 11656 8730
rect 11708 8678 11720 8730
rect 11772 8678 11784 8730
rect 11836 8678 11848 8730
rect 11900 8678 12512 8730
rect 1104 8656 12512 8678
rect 2130 8576 2136 8628
rect 2188 8576 2194 8628
rect 3326 8616 3332 8628
rect 2240 8588 3332 8616
rect 1670 8508 1676 8560
rect 1728 8508 1734 8560
rect 1889 8551 1947 8557
rect 1889 8517 1901 8551
rect 1935 8548 1947 8551
rect 1935 8520 2176 8548
rect 1935 8517 1947 8520
rect 1889 8511 1947 8517
rect 2148 8492 2176 8520
rect 2130 8440 2136 8492
rect 2188 8440 2194 8492
rect 2240 8480 2268 8588
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 3418 8576 3424 8628
rect 3476 8576 3482 8628
rect 3786 8576 3792 8628
rect 3844 8576 3850 8628
rect 3970 8576 3976 8628
rect 4028 8576 4034 8628
rect 4154 8576 4160 8628
rect 4212 8576 4218 8628
rect 5626 8616 5632 8628
rect 5184 8588 5632 8616
rect 2406 8508 2412 8560
rect 2464 8548 2470 8560
rect 2685 8551 2743 8557
rect 2685 8548 2697 8551
rect 2464 8520 2697 8548
rect 2464 8508 2470 8520
rect 2685 8517 2697 8520
rect 2731 8517 2743 8551
rect 3436 8548 3464 8576
rect 3804 8548 3832 8576
rect 5184 8557 5212 8588
rect 5626 8576 5632 8588
rect 5684 8616 5690 8628
rect 7098 8616 7104 8628
rect 5684 8588 7104 8616
rect 5684 8576 5690 8588
rect 5169 8551 5227 8557
rect 2685 8511 2743 8517
rect 3252 8520 3464 8548
rect 3620 8520 3832 8548
rect 4356 8520 4844 8548
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 2240 8452 2329 8480
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 3142 8440 3148 8492
rect 3200 8440 3206 8492
rect 2222 8372 2228 8424
rect 2280 8412 2286 8424
rect 2593 8415 2651 8421
rect 2593 8412 2605 8415
rect 2280 8384 2605 8412
rect 2280 8372 2286 8384
rect 2593 8381 2605 8384
rect 2639 8412 2651 8415
rect 3252 8412 3280 8520
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 3510 8480 3516 8492
rect 3467 8452 3516 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 2639 8384 3280 8412
rect 3329 8415 3387 8421
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3620 8412 3648 8520
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4062 8480 4068 8492
rect 3844 8452 4068 8480
rect 3844 8440 3850 8452
rect 4062 8440 4068 8452
rect 4120 8440 4126 8492
rect 4356 8489 4384 8520
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4430 8440 4436 8492
rect 4488 8440 4494 8492
rect 4709 8483 4767 8489
rect 4709 8449 4721 8483
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 3375 8384 3648 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8344 2099 8347
rect 3344 8344 3372 8375
rect 3970 8372 3976 8424
rect 4028 8412 4034 8424
rect 4724 8412 4752 8443
rect 4028 8384 4752 8412
rect 4028 8372 4034 8384
rect 2087 8316 3372 8344
rect 2087 8313 2099 8316
rect 2041 8307 2099 8313
rect 4522 8304 4528 8356
rect 4580 8344 4586 8356
rect 4617 8347 4675 8353
rect 4617 8344 4629 8347
rect 4580 8316 4629 8344
rect 4580 8304 4586 8316
rect 4617 8313 4629 8316
rect 4663 8313 4675 8347
rect 4816 8344 4844 8520
rect 5169 8517 5181 8551
rect 5215 8517 5227 8551
rect 5169 8511 5227 8517
rect 5258 8508 5264 8560
rect 5316 8548 5322 8560
rect 5316 8520 6132 8548
rect 5316 8508 5322 8520
rect 4890 8440 4896 8492
rect 4948 8440 4954 8492
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8449 5043 8483
rect 4985 8443 5043 8449
rect 5000 8412 5028 8443
rect 5350 8440 5356 8492
rect 5408 8440 5414 8492
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 5629 8415 5687 8421
rect 5629 8412 5641 8415
rect 5000 8384 5641 8412
rect 5629 8381 5641 8384
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 5828 8344 5856 8443
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 6104 8421 6132 8520
rect 6196 8489 6224 8588
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 8018 8576 8024 8628
rect 8076 8576 8082 8628
rect 9582 8576 9588 8628
rect 9640 8616 9646 8628
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 9640 8588 9873 8616
rect 9640 8576 9646 8588
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 9861 8579 9919 8585
rect 11330 8576 11336 8628
rect 11388 8576 11394 8628
rect 11514 8576 11520 8628
rect 11572 8576 11578 8628
rect 8110 8508 8116 8560
rect 8168 8548 8174 8560
rect 9677 8551 9735 8557
rect 8168 8520 8616 8548
rect 8168 8508 8174 8520
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8449 6239 8483
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 6181 8443 6239 8449
rect 6932 8452 8217 8480
rect 6089 8415 6147 8421
rect 6089 8381 6101 8415
rect 6135 8412 6147 8415
rect 6822 8412 6828 8424
rect 6135 8384 6828 8412
rect 6135 8381 6147 8384
rect 6089 8375 6147 8381
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 6362 8344 6368 8356
rect 4816 8316 6368 8344
rect 4617 8307 4675 8313
rect 6362 8304 6368 8316
rect 6420 8344 6426 8356
rect 6932 8344 6960 8452
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8478 8480 8484 8492
rect 8343 8452 8484 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 8588 8489 8616 8520
rect 9677 8517 9689 8551
rect 9723 8548 9735 8551
rect 9723 8520 11836 8548
rect 9723 8517 9735 8520
rect 9677 8511 9735 8517
rect 8573 8483 8631 8489
rect 8573 8449 8585 8483
rect 8619 8480 8631 8483
rect 8619 8452 8708 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 6420 8316 6960 8344
rect 6420 8304 6426 8316
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 8481 8347 8539 8353
rect 8481 8344 8493 8347
rect 7800 8316 8493 8344
rect 7800 8304 7806 8316
rect 8481 8313 8493 8316
rect 8527 8313 8539 8347
rect 8680 8344 8708 8452
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9309 8483 9367 8489
rect 9309 8480 9321 8483
rect 9180 8452 9321 8480
rect 9180 8440 9186 8452
rect 9309 8449 9321 8452
rect 9355 8449 9367 8483
rect 9309 8443 9367 8449
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 9766 8440 9772 8492
rect 9824 8440 9830 8492
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8480 10011 8483
rect 10318 8480 10324 8492
rect 9999 8452 10324 8480
rect 9999 8449 10011 8452
rect 9953 8443 10011 8449
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 10686 8480 10692 8492
rect 10428 8452 10692 8480
rect 9858 8372 9864 8424
rect 9916 8412 9922 8424
rect 10428 8412 10456 8452
rect 10686 8440 10692 8452
rect 10744 8480 10750 8492
rect 11072 8489 11100 8520
rect 11808 8492 11836 8520
rect 10873 8483 10931 8489
rect 10873 8480 10885 8483
rect 10744 8452 10885 8480
rect 10744 8440 10750 8452
rect 10873 8449 10885 8452
rect 10919 8449 10931 8483
rect 10873 8443 10931 8449
rect 11057 8483 11115 8489
rect 11057 8449 11069 8483
rect 11103 8449 11115 8483
rect 11057 8443 11115 8449
rect 11149 8483 11207 8489
rect 11149 8449 11161 8483
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 9916 8384 10456 8412
rect 9916 8372 9922 8384
rect 10778 8372 10784 8424
rect 10836 8412 10842 8424
rect 11164 8412 11192 8443
rect 11790 8440 11796 8492
rect 11848 8440 11854 8492
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 10836 8384 11529 8412
rect 10836 8372 10842 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 11517 8375 11575 8381
rect 8680 8316 9720 8344
rect 8481 8307 8539 8313
rect 1854 8236 1860 8288
rect 1912 8236 1918 8288
rect 2501 8279 2559 8285
rect 2501 8245 2513 8279
rect 2547 8276 2559 8279
rect 2866 8276 2872 8288
rect 2547 8248 2872 8276
rect 2547 8245 2559 8248
rect 2501 8239 2559 8245
rect 2866 8236 2872 8248
rect 2924 8276 2930 8288
rect 3602 8276 3608 8288
rect 2924 8248 3608 8276
rect 2924 8236 2930 8248
rect 3602 8236 3608 8248
rect 3660 8236 3666 8288
rect 3694 8236 3700 8288
rect 3752 8276 3758 8288
rect 5350 8276 5356 8288
rect 3752 8248 5356 8276
rect 3752 8236 3758 8248
rect 5350 8236 5356 8248
rect 5408 8236 5414 8288
rect 5537 8279 5595 8285
rect 5537 8245 5549 8279
rect 5583 8276 5595 8279
rect 5718 8276 5724 8288
rect 5583 8248 5724 8276
rect 5583 8245 5595 8248
rect 5537 8239 5595 8245
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 8294 8276 8300 8288
rect 7248 8248 8300 8276
rect 7248 8236 7254 8248
rect 8294 8236 8300 8248
rect 8352 8236 8358 8288
rect 9692 8276 9720 8316
rect 10318 8304 10324 8356
rect 10376 8344 10382 8356
rect 10965 8347 11023 8353
rect 10965 8344 10977 8347
rect 10376 8316 10977 8344
rect 10376 8304 10382 8316
rect 10965 8313 10977 8316
rect 11011 8344 11023 8347
rect 11330 8344 11336 8356
rect 11011 8316 11336 8344
rect 11011 8313 11023 8316
rect 10965 8307 11023 8313
rect 11330 8304 11336 8316
rect 11388 8344 11394 8356
rect 11701 8347 11759 8353
rect 11701 8344 11713 8347
rect 11388 8316 11713 8344
rect 11388 8304 11394 8316
rect 11701 8313 11713 8316
rect 11747 8313 11759 8347
rect 11701 8307 11759 8313
rect 10502 8276 10508 8288
rect 9692 8248 10508 8276
rect 10502 8236 10508 8248
rect 10560 8236 10566 8288
rect 1104 8186 12512 8208
rect 1104 8134 2376 8186
rect 2428 8134 2440 8186
rect 2492 8134 2504 8186
rect 2556 8134 2568 8186
rect 2620 8134 2632 8186
rect 2684 8134 5228 8186
rect 5280 8134 5292 8186
rect 5344 8134 5356 8186
rect 5408 8134 5420 8186
rect 5472 8134 5484 8186
rect 5536 8134 8080 8186
rect 8132 8134 8144 8186
rect 8196 8134 8208 8186
rect 8260 8134 8272 8186
rect 8324 8134 8336 8186
rect 8388 8134 10932 8186
rect 10984 8134 10996 8186
rect 11048 8134 11060 8186
rect 11112 8134 11124 8186
rect 11176 8134 11188 8186
rect 11240 8134 12512 8186
rect 1104 8112 12512 8134
rect 1302 8032 1308 8084
rect 1360 8072 1366 8084
rect 1857 8075 1915 8081
rect 1857 8072 1869 8075
rect 1360 8044 1869 8072
rect 1360 8032 1366 8044
rect 1857 8041 1869 8044
rect 1903 8041 1915 8075
rect 1857 8035 1915 8041
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2222 8072 2228 8084
rect 2096 8044 2228 8072
rect 2096 8032 2102 8044
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 2593 8075 2651 8081
rect 2593 8041 2605 8075
rect 2639 8072 2651 8075
rect 3510 8072 3516 8084
rect 2639 8044 3516 8072
rect 2639 8041 2651 8044
rect 2593 8035 2651 8041
rect 3510 8032 3516 8044
rect 3568 8032 3574 8084
rect 4430 8032 4436 8084
rect 4488 8072 4494 8084
rect 4801 8075 4859 8081
rect 4801 8072 4813 8075
rect 4488 8044 4813 8072
rect 4488 8032 4494 8044
rect 4801 8041 4813 8044
rect 4847 8041 4859 8075
rect 4801 8035 4859 8041
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 5902 8072 5908 8084
rect 5491 8044 5908 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 7929 8075 7987 8081
rect 7929 8041 7941 8075
rect 7975 8072 7987 8075
rect 9490 8072 9496 8084
rect 7975 8044 9496 8072
rect 7975 8041 7987 8044
rect 7929 8035 7987 8041
rect 9490 8032 9496 8044
rect 9548 8032 9554 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10836 8044 10885 8072
rect 10836 8032 10842 8044
rect 10873 8041 10885 8044
rect 10919 8041 10931 8075
rect 10873 8035 10931 8041
rect 1486 7964 1492 8016
rect 1544 7964 1550 8016
rect 1670 7964 1676 8016
rect 1728 8004 1734 8016
rect 2498 8004 2504 8016
rect 1728 7976 2504 8004
rect 1728 7964 1734 7976
rect 2498 7964 2504 7976
rect 2556 7964 2562 8016
rect 2777 8007 2835 8013
rect 2777 7973 2789 8007
rect 2823 8004 2835 8007
rect 2866 8004 2872 8016
rect 2823 7976 2872 8004
rect 2823 7973 2835 7976
rect 2777 7967 2835 7973
rect 2866 7964 2872 7976
rect 2924 7964 2930 8016
rect 10962 7964 10968 8016
rect 11020 7964 11026 8016
rect 4982 7936 4988 7948
rect 1688 7908 4988 7936
rect 1688 7877 1716 7908
rect 4982 7896 4988 7908
rect 5040 7896 5046 7948
rect 6546 7896 6552 7948
rect 6604 7936 6610 7948
rect 7469 7939 7527 7945
rect 7469 7936 7481 7939
rect 6604 7908 7481 7936
rect 6604 7896 6610 7908
rect 7469 7905 7481 7908
rect 7515 7905 7527 7939
rect 7469 7899 7527 7905
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 2038 7828 2044 7880
rect 2096 7828 2102 7880
rect 2130 7828 2136 7880
rect 2188 7868 2194 7880
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 2188 7840 2329 7868
rect 2188 7828 2194 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 2593 7871 2651 7877
rect 2593 7868 2605 7871
rect 2556 7840 2605 7868
rect 2556 7828 2562 7840
rect 2593 7837 2605 7840
rect 2639 7837 2651 7871
rect 2593 7831 2651 7837
rect 2682 7828 2688 7880
rect 2740 7828 2746 7880
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 3878 7868 3884 7880
rect 2915 7840 3884 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 1854 7760 1860 7812
rect 1912 7800 1918 7812
rect 2409 7803 2467 7809
rect 2409 7800 2421 7803
rect 1912 7772 2421 7800
rect 1912 7760 1918 7772
rect 2409 7769 2421 7772
rect 2455 7769 2467 7803
rect 2409 7763 2467 7769
rect 2424 7732 2452 7763
rect 2884 7744 2912 7831
rect 3878 7828 3884 7840
rect 3936 7828 3942 7880
rect 4522 7828 4528 7880
rect 4580 7828 4586 7880
rect 5074 7828 5080 7880
rect 5132 7868 5138 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 5132 7840 5181 7868
rect 5132 7828 5138 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5626 7868 5632 7880
rect 5307 7840 5632 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7561 7871 7619 7877
rect 7561 7868 7573 7871
rect 7156 7840 7573 7868
rect 7156 7828 7162 7840
rect 7561 7837 7573 7840
rect 7607 7868 7619 7871
rect 8110 7868 8116 7880
rect 7607 7840 8116 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 8110 7828 8116 7840
rect 8168 7828 8174 7880
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 3970 7760 3976 7812
rect 4028 7800 4034 7812
rect 4617 7803 4675 7809
rect 4617 7800 4629 7803
rect 4028 7772 4629 7800
rect 4028 7760 4034 7772
rect 4617 7769 4629 7772
rect 4663 7769 4675 7803
rect 4617 7763 4675 7769
rect 4801 7803 4859 7809
rect 4801 7769 4813 7803
rect 4847 7800 4859 7803
rect 5445 7803 5503 7809
rect 5445 7800 5457 7803
rect 4847 7772 5457 7800
rect 4847 7769 4859 7772
rect 4801 7763 4859 7769
rect 5092 7744 5120 7772
rect 5445 7769 5457 7772
rect 5491 7769 5503 7803
rect 10336 7800 10364 7831
rect 10410 7828 10416 7880
rect 10468 7828 10474 7880
rect 11790 7828 11796 7880
rect 11848 7828 11854 7880
rect 10502 7800 10508 7812
rect 10336 7772 10508 7800
rect 5445 7763 5503 7769
rect 10502 7760 10508 7772
rect 10560 7760 10566 7812
rect 10597 7803 10655 7809
rect 10597 7769 10609 7803
rect 10643 7800 10655 7803
rect 11333 7803 11391 7809
rect 11333 7800 11345 7803
rect 10643 7772 11345 7800
rect 10643 7769 10655 7772
rect 10597 7763 10655 7769
rect 11333 7769 11345 7772
rect 11379 7800 11391 7803
rect 11609 7803 11667 7809
rect 11609 7800 11621 7803
rect 11379 7772 11621 7800
rect 11379 7769 11391 7772
rect 11333 7763 11391 7769
rect 11609 7769 11621 7772
rect 11655 7769 11667 7803
rect 11609 7763 11667 7769
rect 2866 7732 2872 7744
rect 2424 7704 2872 7732
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 5074 7692 5080 7744
rect 5132 7692 5138 7744
rect 7193 7735 7251 7741
rect 7193 7701 7205 7735
rect 7239 7732 7251 7735
rect 7926 7732 7932 7744
rect 7239 7704 7932 7732
rect 7239 7701 7251 7704
rect 7193 7695 7251 7701
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 11422 7692 11428 7744
rect 11480 7692 11486 7744
rect 1104 7642 12512 7664
rect 1104 7590 3036 7642
rect 3088 7590 3100 7642
rect 3152 7590 3164 7642
rect 3216 7590 3228 7642
rect 3280 7590 3292 7642
rect 3344 7590 5888 7642
rect 5940 7590 5952 7642
rect 6004 7590 6016 7642
rect 6068 7590 6080 7642
rect 6132 7590 6144 7642
rect 6196 7590 8740 7642
rect 8792 7590 8804 7642
rect 8856 7590 8868 7642
rect 8920 7590 8932 7642
rect 8984 7590 8996 7642
rect 9048 7590 11592 7642
rect 11644 7590 11656 7642
rect 11708 7590 11720 7642
rect 11772 7590 11784 7642
rect 11836 7590 11848 7642
rect 11900 7590 12512 7642
rect 1104 7568 12512 7590
rect 1949 7531 2007 7537
rect 1949 7497 1961 7531
rect 1995 7528 2007 7531
rect 1995 7500 5028 7528
rect 1995 7497 2007 7500
rect 1949 7491 2007 7497
rect 934 7420 940 7472
rect 992 7460 998 7472
rect 2317 7463 2375 7469
rect 992 7432 1808 7460
rect 992 7420 998 7432
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 1780 7401 1808 7432
rect 2317 7429 2329 7463
rect 2363 7460 2375 7463
rect 2866 7460 2872 7472
rect 2363 7432 2872 7460
rect 2363 7429 2375 7432
rect 2317 7423 2375 7429
rect 2866 7420 2872 7432
rect 2924 7420 2930 7472
rect 3053 7463 3111 7469
rect 3053 7429 3065 7463
rect 3099 7460 3111 7463
rect 3970 7460 3976 7472
rect 3099 7432 3976 7460
rect 3099 7429 3111 7432
rect 3053 7423 3111 7429
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 5000 7469 5028 7500
rect 6546 7488 6552 7540
rect 6604 7488 6610 7540
rect 7745 7531 7803 7537
rect 7745 7497 7757 7531
rect 7791 7528 7803 7531
rect 10410 7528 10416 7540
rect 7791 7500 10416 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 10336 7469 10364 7500
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 11514 7528 11520 7540
rect 10612 7500 11520 7528
rect 4985 7463 5043 7469
rect 4985 7429 4997 7463
rect 5031 7460 5043 7463
rect 10321 7463 10379 7469
rect 5031 7432 5488 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 1946 7352 1952 7404
rect 2004 7392 2010 7404
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 2004 7364 2513 7392
rect 2004 7352 2010 7364
rect 2501 7361 2513 7364
rect 2547 7392 2559 7395
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2547 7364 2789 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 2682 7284 2688 7336
rect 2740 7284 2746 7336
rect 2792 7324 2820 7355
rect 3326 7352 3332 7404
rect 3384 7352 3390 7404
rect 3786 7352 3792 7404
rect 3844 7392 3850 7404
rect 5460 7401 5488 7432
rect 10321 7429 10333 7463
rect 10367 7429 10379 7463
rect 10321 7423 10379 7429
rect 10502 7420 10508 7472
rect 10560 7420 10566 7472
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 3844 7364 5181 7392
rect 3844 7352 3850 7364
rect 5169 7361 5181 7364
rect 5215 7361 5227 7395
rect 5169 7355 5227 7361
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 3344 7324 3372 7352
rect 2792 7296 3372 7324
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7324 5411 7327
rect 6380 7324 6408 7355
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 6730 7392 6736 7404
rect 6604 7364 6736 7392
rect 6604 7352 6610 7364
rect 6730 7352 6736 7364
rect 6788 7392 6794 7404
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 6788 7364 6929 7392
rect 6788 7352 6794 7364
rect 6917 7361 6929 7364
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 5399 7296 6408 7324
rect 5399 7293 5411 7296
rect 5353 7287 5411 7293
rect 2130 7216 2136 7268
rect 2188 7256 2194 7268
rect 2700 7256 2728 7284
rect 3237 7259 3295 7265
rect 3237 7256 3249 7259
rect 2188 7228 3249 7256
rect 2188 7216 2194 7228
rect 3237 7225 3249 7228
rect 3283 7225 3295 7259
rect 3237 7219 3295 7225
rect 3878 7216 3884 7268
rect 3936 7256 3942 7268
rect 5629 7259 5687 7265
rect 5629 7256 5641 7259
rect 3936 7228 5641 7256
rect 3936 7216 3942 7228
rect 5629 7225 5641 7228
rect 5675 7225 5687 7259
rect 6380 7256 6408 7296
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 7006 7324 7012 7336
rect 6687 7296 7012 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 7147 7296 7297 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7285 7293 7297 7296
rect 7331 7293 7343 7327
rect 7392 7324 7420 7355
rect 7926 7352 7932 7404
rect 7984 7352 7990 7404
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 8076 7364 8217 7392
rect 8076 7352 8082 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 10134 7352 10140 7404
rect 10192 7392 10198 7404
rect 10612 7392 10640 7500
rect 11514 7488 11520 7500
rect 11572 7528 11578 7540
rect 11701 7531 11759 7537
rect 11701 7528 11713 7531
rect 11572 7500 11713 7528
rect 11572 7488 11578 7500
rect 11701 7497 11713 7500
rect 11747 7497 11759 7531
rect 11701 7491 11759 7497
rect 10192 7364 10640 7392
rect 10192 7352 10198 7364
rect 10686 7352 10692 7404
rect 10744 7392 10750 7404
rect 10962 7392 10968 7404
rect 10744 7364 10968 7392
rect 10744 7352 10750 7364
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7392 11207 7395
rect 11422 7392 11428 7404
rect 11195 7364 11428 7392
rect 11195 7361 11207 7364
rect 11149 7355 11207 7361
rect 11422 7352 11428 7364
rect 11480 7352 11486 7404
rect 11514 7352 11520 7404
rect 11572 7352 11578 7404
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 11974 7392 11980 7404
rect 11839 7364 11980 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 7834 7324 7840 7336
rect 7392 7296 7840 7324
rect 7285 7287 7343 7293
rect 7834 7284 7840 7296
rect 7892 7324 7898 7336
rect 8036 7324 8064 7352
rect 7892 7296 8064 7324
rect 7892 7284 7898 7296
rect 8110 7284 8116 7336
rect 8168 7284 8174 7336
rect 11241 7327 11299 7333
rect 11241 7293 11253 7327
rect 11287 7324 11299 7327
rect 11330 7324 11336 7336
rect 11287 7296 11336 7324
rect 11287 7293 11299 7296
rect 11241 7287 11299 7293
rect 11330 7284 11336 7296
rect 11388 7284 11394 7336
rect 6733 7259 6791 7265
rect 6733 7256 6745 7259
rect 6380 7228 6745 7256
rect 5629 7219 5687 7225
rect 6733 7225 6745 7228
rect 6779 7256 6791 7259
rect 7466 7256 7472 7268
rect 6779 7228 7472 7256
rect 6779 7225 6791 7228
rect 6733 7219 6791 7225
rect 7466 7216 7472 7228
rect 7524 7256 7530 7268
rect 8021 7259 8079 7265
rect 8021 7256 8033 7259
rect 7524 7228 8033 7256
rect 7524 7216 7530 7228
rect 8021 7225 8033 7228
rect 8067 7225 8079 7259
rect 8021 7219 8079 7225
rect 10870 7216 10876 7268
rect 10928 7256 10934 7268
rect 11517 7259 11575 7265
rect 11517 7256 11529 7259
rect 10928 7228 11529 7256
rect 10928 7216 10934 7228
rect 11517 7225 11529 7228
rect 11563 7225 11575 7259
rect 11517 7219 11575 7225
rect 1486 7148 1492 7200
rect 1544 7148 1550 7200
rect 2222 7148 2228 7200
rect 2280 7188 2286 7200
rect 2685 7191 2743 7197
rect 2685 7188 2697 7191
rect 2280 7160 2697 7188
rect 2280 7148 2286 7160
rect 2685 7157 2697 7160
rect 2731 7157 2743 7191
rect 2685 7151 2743 7157
rect 2774 7148 2780 7200
rect 2832 7148 2838 7200
rect 8389 7191 8447 7197
rect 8389 7157 8401 7191
rect 8435 7188 8447 7191
rect 8478 7188 8484 7200
rect 8435 7160 8484 7188
rect 8435 7157 8447 7160
rect 8389 7151 8447 7157
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 9950 7148 9956 7200
rect 10008 7188 10014 7200
rect 10781 7191 10839 7197
rect 10781 7188 10793 7191
rect 10008 7160 10793 7188
rect 10008 7148 10014 7160
rect 10781 7157 10793 7160
rect 10827 7157 10839 7191
rect 10781 7151 10839 7157
rect 1104 7098 12512 7120
rect 1104 7046 2376 7098
rect 2428 7046 2440 7098
rect 2492 7046 2504 7098
rect 2556 7046 2568 7098
rect 2620 7046 2632 7098
rect 2684 7046 5228 7098
rect 5280 7046 5292 7098
rect 5344 7046 5356 7098
rect 5408 7046 5420 7098
rect 5472 7046 5484 7098
rect 5536 7046 8080 7098
rect 8132 7046 8144 7098
rect 8196 7046 8208 7098
rect 8260 7046 8272 7098
rect 8324 7046 8336 7098
rect 8388 7046 10932 7098
rect 10984 7046 10996 7098
rect 11048 7046 11060 7098
rect 11112 7046 11124 7098
rect 11176 7046 11188 7098
rect 11240 7046 12512 7098
rect 1104 7024 12512 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 2133 6987 2191 6993
rect 2133 6984 2145 6987
rect 1728 6956 2145 6984
rect 1728 6944 1734 6956
rect 2133 6953 2145 6956
rect 2179 6953 2191 6987
rect 2133 6947 2191 6953
rect 7466 6944 7472 6996
rect 7524 6944 7530 6996
rect 5350 6916 5356 6928
rect 2528 6888 5356 6916
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 2528 6780 2556 6888
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 7006 6876 7012 6928
rect 7064 6916 7070 6928
rect 7561 6919 7619 6925
rect 7561 6916 7573 6919
rect 7064 6888 7573 6916
rect 7064 6876 7070 6888
rect 7561 6885 7573 6888
rect 7607 6885 7619 6919
rect 7561 6879 7619 6885
rect 10042 6876 10048 6928
rect 10100 6916 10106 6928
rect 11974 6916 11980 6928
rect 10100 6888 11980 6916
rect 10100 6876 10106 6888
rect 11974 6876 11980 6888
rect 12032 6876 12038 6928
rect 2866 6808 2872 6860
rect 2924 6848 2930 6860
rect 7926 6848 7932 6860
rect 2924 6820 3464 6848
rect 2924 6808 2930 6820
rect 2363 6752 2556 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2648 6752 2697 6780
rect 2648 6740 2654 6752
rect 2685 6749 2697 6752
rect 2731 6749 2743 6783
rect 2685 6743 2743 6749
rect 3053 6783 3111 6789
rect 3053 6749 3065 6783
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 3145 6783 3203 6789
rect 3145 6749 3157 6783
rect 3191 6749 3203 6783
rect 3145 6743 3203 6749
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3326 6780 3332 6792
rect 3283 6752 3332 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 2130 6672 2136 6724
rect 2188 6712 2194 6724
rect 2409 6715 2467 6721
rect 2409 6712 2421 6715
rect 2188 6684 2421 6712
rect 2188 6672 2194 6684
rect 2409 6681 2421 6684
rect 2455 6681 2467 6715
rect 2409 6675 2467 6681
rect 2501 6715 2559 6721
rect 2501 6681 2513 6715
rect 2547 6681 2559 6715
rect 2501 6675 2559 6681
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 2516 6644 2544 6675
rect 2280 6616 2544 6644
rect 2777 6647 2835 6653
rect 2280 6604 2286 6616
rect 2777 6613 2789 6647
rect 2823 6644 2835 6647
rect 2958 6644 2964 6656
rect 2823 6616 2964 6644
rect 2823 6613 2835 6616
rect 2777 6607 2835 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3068 6644 3096 6743
rect 3160 6712 3188 6743
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3436 6789 3464 6820
rect 7392 6820 7932 6848
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 7392 6789 7420 6820
rect 7926 6808 7932 6820
rect 7984 6808 7990 6860
rect 8389 6851 8447 6857
rect 8389 6848 8401 6851
rect 8220 6820 8401 6848
rect 5169 6783 5227 6789
rect 5169 6780 5181 6783
rect 4948 6752 5181 6780
rect 4948 6740 4954 6752
rect 5169 6749 5181 6752
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7653 6783 7711 6789
rect 7653 6749 7665 6783
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 3694 6712 3700 6724
rect 3160 6684 3700 6712
rect 3694 6672 3700 6684
rect 3752 6712 3758 6724
rect 7190 6712 7196 6724
rect 3752 6684 7196 6712
rect 3752 6672 3758 6684
rect 5184 6656 5212 6684
rect 7190 6672 7196 6684
rect 7248 6712 7254 6724
rect 7668 6712 7696 6743
rect 7834 6740 7840 6792
rect 7892 6740 7898 6792
rect 8220 6712 8248 6820
rect 8389 6817 8401 6820
rect 8435 6848 8447 6851
rect 10502 6848 10508 6860
rect 8435 6820 9260 6848
rect 8435 6817 8447 6820
rect 8389 6811 8447 6817
rect 8297 6783 8355 6789
rect 8297 6749 8309 6783
rect 8343 6780 8355 6783
rect 8478 6780 8484 6792
rect 8343 6752 8484 6780
rect 8343 6749 8355 6752
rect 8297 6743 8355 6749
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 9232 6724 9260 6820
rect 9784 6820 10508 6848
rect 9784 6789 9812 6820
rect 10502 6808 10508 6820
rect 10560 6848 10566 6860
rect 10597 6851 10655 6857
rect 10597 6848 10609 6851
rect 10560 6820 10609 6848
rect 10560 6808 10566 6820
rect 10597 6817 10609 6820
rect 10643 6817 10655 6851
rect 11422 6848 11428 6860
rect 10597 6811 10655 6817
rect 11072 6820 11428 6848
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 10042 6740 10048 6792
rect 10100 6740 10106 6792
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 11072 6789 11100 6820
rect 11422 6808 11428 6820
rect 11480 6808 11486 6860
rect 12158 6808 12164 6860
rect 12216 6808 12222 6860
rect 11057 6783 11115 6789
rect 11057 6749 11069 6783
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6780 11299 6783
rect 11330 6780 11336 6792
rect 11287 6752 11336 6780
rect 11287 6749 11299 6752
rect 11241 6743 11299 6749
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 11885 6783 11943 6789
rect 11885 6749 11897 6783
rect 11931 6749 11943 6783
rect 11885 6743 11943 6749
rect 7248 6684 7604 6712
rect 7668 6684 8248 6712
rect 7248 6672 7254 6684
rect 3786 6644 3792 6656
rect 3068 6616 3792 6644
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 5166 6604 5172 6656
rect 5224 6604 5230 6656
rect 5350 6604 5356 6656
rect 5408 6644 5414 6656
rect 6270 6644 6276 6656
rect 5408 6616 6276 6644
rect 5408 6604 5414 6616
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 7101 6647 7159 6653
rect 7101 6613 7113 6647
rect 7147 6644 7159 6647
rect 7466 6644 7472 6656
rect 7147 6616 7472 6644
rect 7147 6613 7159 6616
rect 7101 6607 7159 6613
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 7576 6644 7604 6684
rect 9214 6672 9220 6724
rect 9272 6712 9278 6724
rect 11900 6712 11928 6743
rect 9272 6684 11928 6712
rect 9272 6672 9278 6684
rect 8478 6644 8484 6656
rect 7576 6616 8484 6644
rect 8478 6604 8484 6616
rect 8536 6604 8542 6656
rect 8665 6647 8723 6653
rect 8665 6613 8677 6647
rect 8711 6644 8723 6647
rect 9490 6644 9496 6656
rect 8711 6616 9496 6644
rect 8711 6613 8723 6616
rect 8665 6607 8723 6613
rect 9490 6604 9496 6616
rect 9548 6604 9554 6656
rect 9585 6647 9643 6653
rect 9585 6613 9597 6647
rect 9631 6644 9643 6647
rect 10962 6644 10968 6656
rect 9631 6616 10968 6644
rect 9631 6613 9643 6616
rect 9585 6607 9643 6613
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 1104 6554 12512 6576
rect 1104 6502 3036 6554
rect 3088 6502 3100 6554
rect 3152 6502 3164 6554
rect 3216 6502 3228 6554
rect 3280 6502 3292 6554
rect 3344 6502 5888 6554
rect 5940 6502 5952 6554
rect 6004 6502 6016 6554
rect 6068 6502 6080 6554
rect 6132 6502 6144 6554
rect 6196 6502 8740 6554
rect 8792 6502 8804 6554
rect 8856 6502 8868 6554
rect 8920 6502 8932 6554
rect 8984 6502 8996 6554
rect 9048 6502 11592 6554
rect 11644 6502 11656 6554
rect 11708 6502 11720 6554
rect 11772 6502 11784 6554
rect 11836 6502 11848 6554
rect 11900 6502 12512 6554
rect 1104 6480 12512 6502
rect 2590 6400 2596 6452
rect 2648 6400 2654 6452
rect 3513 6443 3571 6449
rect 3513 6409 3525 6443
rect 3559 6440 3571 6443
rect 4890 6440 4896 6452
rect 3559 6412 4896 6440
rect 3559 6409 3571 6412
rect 3513 6403 3571 6409
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 7098 6440 7104 6452
rect 5368 6412 7104 6440
rect 2958 6332 2964 6384
rect 3016 6372 3022 6384
rect 4908 6372 4936 6400
rect 5368 6372 5396 6412
rect 7098 6400 7104 6412
rect 7156 6440 7162 6452
rect 7374 6440 7380 6452
rect 7156 6412 7380 6440
rect 7156 6400 7162 6412
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 8665 6443 8723 6449
rect 8128 6412 8616 6440
rect 3016 6344 3096 6372
rect 3016 6332 3022 6344
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1489 6307 1547 6313
rect 1489 6304 1501 6307
rect 900 6276 1501 6304
rect 900 6264 906 6276
rect 1489 6273 1501 6276
rect 1535 6273 1547 6307
rect 1489 6267 1547 6273
rect 2774 6264 2780 6316
rect 2832 6264 2838 6316
rect 3068 6313 3096 6344
rect 3436 6344 3832 6372
rect 4908 6344 5396 6372
rect 3436 6313 3464 6344
rect 3804 6313 3832 6344
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3513 6307 3571 6313
rect 3513 6273 3525 6307
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6273 3847 6307
rect 3789 6267 3847 6273
rect 2866 6196 2872 6248
rect 2924 6196 2930 6248
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3142 6236 3148 6248
rect 3007 6208 3148 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 3142 6196 3148 6208
rect 3200 6236 3206 6248
rect 3436 6236 3464 6267
rect 3200 6208 3464 6236
rect 3200 6196 3206 6208
rect 3528 6168 3556 6267
rect 4062 6264 4068 6316
rect 4120 6264 4126 6316
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 4764 6276 5089 6304
rect 4764 6264 4770 6276
rect 5077 6273 5089 6276
rect 5123 6273 5135 6307
rect 5077 6267 5135 6273
rect 5166 6264 5172 6316
rect 5224 6264 5230 6316
rect 5368 6304 5396 6344
rect 6362 6332 6368 6384
rect 6420 6372 6426 6384
rect 8128 6372 8156 6412
rect 6420 6344 8156 6372
rect 8220 6344 8432 6372
rect 6420 6332 6426 6344
rect 5435 6307 5493 6313
rect 5435 6304 5447 6307
rect 5368 6276 5447 6304
rect 5435 6273 5447 6276
rect 5481 6273 5493 6307
rect 5435 6267 5493 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 5721 6307 5779 6313
rect 5721 6273 5733 6307
rect 5767 6273 5779 6307
rect 5721 6267 5779 6273
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 3436 6140 3556 6168
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6100 1823 6103
rect 2774 6100 2780 6112
rect 1811 6072 2780 6100
rect 1811 6069 1823 6072
rect 1765 6063 1823 6069
rect 2774 6060 2780 6072
rect 2832 6100 2838 6112
rect 3436 6100 3464 6140
rect 3786 6128 3792 6180
rect 3844 6128 3850 6180
rect 4908 6168 4936 6199
rect 4982 6196 4988 6248
rect 5040 6196 5046 6248
rect 5353 6239 5411 6245
rect 5353 6205 5365 6239
rect 5399 6236 5411 6239
rect 5552 6236 5580 6267
rect 5399 6208 5580 6236
rect 5736 6236 5764 6267
rect 5810 6264 5816 6316
rect 5868 6264 5874 6316
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7156 6276 8033 6304
rect 7156 6264 7162 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8021 6267 8079 6273
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 7374 6236 7380 6248
rect 5736 6208 7380 6236
rect 5399 6205 5411 6208
rect 5353 6199 5411 6205
rect 5442 6168 5448 6180
rect 4908 6140 5448 6168
rect 5442 6128 5448 6140
rect 5500 6128 5506 6180
rect 5736 6168 5764 6208
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 5552 6140 5764 6168
rect 2832 6072 3464 6100
rect 3804 6100 3832 6128
rect 4798 6100 4804 6112
rect 3804 6072 4804 6100
rect 2832 6060 2838 6072
rect 4798 6060 4804 6072
rect 4856 6100 4862 6112
rect 5552 6100 5580 6140
rect 4856 6072 5580 6100
rect 4856 6060 4862 6072
rect 5626 6060 5632 6112
rect 5684 6100 5690 6112
rect 5997 6103 6055 6109
rect 5997 6100 6009 6103
rect 5684 6072 6009 6100
rect 5684 6060 5690 6072
rect 5997 6069 6009 6072
rect 6043 6069 6055 6103
rect 8128 6100 8156 6267
rect 8220 6168 8248 6344
rect 8404 6313 8432 6344
rect 8297 6307 8355 6313
rect 8297 6273 8309 6307
rect 8343 6273 8355 6307
rect 8297 6267 8355 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 8312 6236 8340 6267
rect 8478 6264 8484 6316
rect 8536 6264 8542 6316
rect 8588 6304 8616 6412
rect 8665 6409 8677 6443
rect 8711 6440 8723 6443
rect 8711 6412 10916 6440
rect 8711 6409 8723 6412
rect 8665 6403 8723 6409
rect 9490 6332 9496 6384
rect 9548 6372 9554 6384
rect 9548 6344 9812 6372
rect 9548 6332 9554 6344
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8588 6276 8953 6304
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 9784 6313 9812 6344
rect 9968 6344 10640 6372
rect 9968 6313 9996 6344
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6304 9367 6307
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 9355 6276 9597 6304
rect 9355 6273 9367 6276
rect 9309 6267 9367 6273
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6304 9827 6307
rect 9861 6307 9919 6313
rect 9861 6304 9873 6307
rect 9815 6276 9873 6304
rect 9815 6273 9827 6276
rect 9769 6267 9827 6273
rect 9861 6273 9873 6276
rect 9907 6273 9919 6307
rect 9861 6267 9919 6273
rect 9953 6307 10011 6313
rect 9953 6273 9965 6307
rect 9999 6273 10011 6307
rect 9953 6267 10011 6273
rect 8570 6236 8576 6248
rect 8312 6208 8576 6236
rect 8570 6196 8576 6208
rect 8628 6236 8634 6248
rect 9324 6236 9352 6267
rect 8628 6208 9352 6236
rect 9600 6236 9628 6267
rect 9968 6236 9996 6267
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10612 6313 10640 6344
rect 10778 6332 10784 6384
rect 10836 6332 10842 6384
rect 10888 6372 10916 6412
rect 10962 6400 10968 6452
rect 11020 6400 11026 6452
rect 11333 6443 11391 6449
rect 11333 6409 11345 6443
rect 11379 6440 11391 6443
rect 11514 6440 11520 6452
rect 11379 6412 11520 6440
rect 11379 6409 11391 6412
rect 11333 6403 11391 6409
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 10888 6344 11192 6372
rect 11164 6313 11192 6344
rect 11974 6332 11980 6384
rect 12032 6332 12038 6384
rect 10505 6307 10563 6313
rect 10505 6304 10517 6307
rect 10284 6276 10517 6304
rect 10284 6264 10290 6276
rect 10505 6273 10517 6276
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 10873 6307 10931 6313
rect 10643 6276 10732 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 9600 6208 9996 6236
rect 8628 6196 8634 6208
rect 10410 6196 10416 6248
rect 10468 6196 10474 6248
rect 9214 6168 9220 6180
rect 8220 6140 9220 6168
rect 9214 6128 9220 6140
rect 9272 6128 9278 6180
rect 10704 6168 10732 6276
rect 10873 6273 10885 6307
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6273 11207 6307
rect 11149 6267 11207 6273
rect 10888 6236 10916 6267
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 10888 6208 11529 6236
rect 11517 6205 11529 6208
rect 11563 6205 11575 6239
rect 11517 6199 11575 6205
rect 11330 6168 11336 6180
rect 10704 6140 11336 6168
rect 11330 6128 11336 6140
rect 11388 6128 11394 6180
rect 11606 6128 11612 6180
rect 11664 6128 11670 6180
rect 8757 6103 8815 6109
rect 8757 6100 8769 6103
rect 8128 6072 8769 6100
rect 5997 6063 6055 6069
rect 8757 6069 8769 6072
rect 8803 6069 8815 6103
rect 8757 6063 8815 6069
rect 9766 6060 9772 6112
rect 9824 6060 9830 6112
rect 10781 6103 10839 6109
rect 10781 6069 10793 6103
rect 10827 6100 10839 6103
rect 11422 6100 11428 6112
rect 10827 6072 11428 6100
rect 10827 6069 10839 6072
rect 10781 6063 10839 6069
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 1104 6010 12512 6032
rect 1104 5958 2376 6010
rect 2428 5958 2440 6010
rect 2492 5958 2504 6010
rect 2556 5958 2568 6010
rect 2620 5958 2632 6010
rect 2684 5958 5228 6010
rect 5280 5958 5292 6010
rect 5344 5958 5356 6010
rect 5408 5958 5420 6010
rect 5472 5958 5484 6010
rect 5536 5958 8080 6010
rect 8132 5958 8144 6010
rect 8196 5958 8208 6010
rect 8260 5958 8272 6010
rect 8324 5958 8336 6010
rect 8388 5958 10932 6010
rect 10984 5958 10996 6010
rect 11048 5958 11060 6010
rect 11112 5958 11124 6010
rect 11176 5958 11188 6010
rect 11240 5958 12512 6010
rect 1104 5936 12512 5958
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 3142 5896 3148 5908
rect 2455 5868 3148 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3329 5899 3387 5905
rect 3329 5865 3341 5899
rect 3375 5896 3387 5899
rect 3418 5896 3424 5908
rect 3375 5868 3424 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 3418 5856 3424 5868
rect 3476 5856 3482 5908
rect 4706 5856 4712 5908
rect 4764 5896 4770 5908
rect 4764 5868 5212 5896
rect 4764 5856 4770 5868
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 3694 5828 3700 5840
rect 2823 5800 3700 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 3694 5788 3700 5800
rect 3752 5788 3758 5840
rect 4985 5831 5043 5837
rect 4985 5797 4997 5831
rect 5031 5797 5043 5831
rect 5184 5828 5212 5868
rect 5626 5856 5632 5908
rect 5684 5856 5690 5908
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 5776 5868 5825 5896
rect 5776 5856 5782 5868
rect 5813 5865 5825 5868
rect 5859 5865 5871 5899
rect 5813 5859 5871 5865
rect 5994 5856 6000 5908
rect 6052 5896 6058 5908
rect 6362 5896 6368 5908
rect 6052 5868 6368 5896
rect 6052 5856 6058 5868
rect 6362 5856 6368 5868
rect 6420 5856 6426 5908
rect 8481 5899 8539 5905
rect 8481 5865 8493 5899
rect 8527 5896 8539 5899
rect 9030 5896 9036 5908
rect 8527 5868 9036 5896
rect 8527 5865 8539 5868
rect 8481 5859 8539 5865
rect 9030 5856 9036 5868
rect 9088 5856 9094 5908
rect 10502 5856 10508 5908
rect 10560 5896 10566 5908
rect 11057 5899 11115 5905
rect 11057 5896 11069 5899
rect 10560 5868 11069 5896
rect 10560 5856 10566 5868
rect 11057 5865 11069 5868
rect 11103 5865 11115 5899
rect 11057 5859 11115 5865
rect 6273 5831 6331 5837
rect 6273 5828 6285 5831
rect 5184 5800 6285 5828
rect 4985 5791 5043 5797
rect 6273 5797 6285 5800
rect 6319 5797 6331 5831
rect 6273 5791 6331 5797
rect 3510 5760 3516 5772
rect 2056 5732 3516 5760
rect 2056 5701 2084 5732
rect 3510 5720 3516 5732
rect 3568 5760 3574 5772
rect 4341 5763 4399 5769
rect 4341 5760 4353 5763
rect 3568 5732 3832 5760
rect 3568 5720 3574 5732
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 2041 5695 2099 5701
rect 2041 5692 2053 5695
rect 1719 5664 2053 5692
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 2041 5661 2053 5664
rect 2087 5661 2099 5695
rect 2041 5655 2099 5661
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2682 5692 2688 5704
rect 2639 5664 2688 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 1486 5584 1492 5636
rect 1544 5584 1550 5636
rect 2222 5584 2228 5636
rect 2280 5584 2286 5636
rect 2608 5624 2636 5655
rect 2682 5652 2688 5664
rect 2740 5652 2746 5704
rect 2777 5695 2835 5701
rect 2777 5661 2789 5695
rect 2823 5692 2835 5695
rect 2866 5692 2872 5704
rect 2823 5664 2872 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 2866 5652 2872 5664
rect 2924 5652 2930 5704
rect 3804 5701 3832 5732
rect 3988 5732 4353 5760
rect 3988 5704 4016 5732
rect 4341 5729 4353 5732
rect 4387 5729 4399 5763
rect 5000 5760 5028 5791
rect 10410 5788 10416 5840
rect 10468 5828 10474 5840
rect 10468 5800 11284 5828
rect 10468 5788 10474 5800
rect 9214 5760 9220 5772
rect 5000 5732 6132 5760
rect 4341 5723 4399 5729
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 4120 5664 4261 5692
rect 4120 5652 4126 5664
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4430 5652 4436 5704
rect 4488 5652 4494 5704
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 4890 5692 4896 5704
rect 4847 5664 4896 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 4890 5652 4896 5664
rect 4948 5692 4954 5704
rect 5202 5695 5260 5701
rect 5202 5692 5214 5695
rect 4948 5664 5214 5692
rect 4948 5652 4954 5664
rect 5202 5661 5214 5664
rect 5248 5692 5260 5695
rect 5721 5695 5779 5701
rect 5248 5664 5672 5692
rect 5248 5661 5260 5664
rect 5202 5655 5260 5661
rect 2961 5627 3019 5633
rect 2961 5624 2973 5627
rect 2608 5596 2973 5624
rect 2961 5593 2973 5596
rect 3007 5593 3019 5627
rect 2961 5587 3019 5593
rect 4154 5584 4160 5636
rect 4212 5584 4218 5636
rect 4522 5584 4528 5636
rect 4580 5624 4586 5636
rect 4985 5627 5043 5633
rect 4580 5596 4936 5624
rect 4580 5584 4586 5596
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3145 5559 3203 5565
rect 3145 5556 3157 5559
rect 2924 5528 3157 5556
rect 2924 5516 2930 5528
rect 3145 5525 3157 5528
rect 3191 5525 3203 5559
rect 3145 5519 3203 5525
rect 3418 5516 3424 5568
rect 3476 5556 3482 5568
rect 4338 5556 4344 5568
rect 3476 5528 4344 5556
rect 3476 5516 3482 5528
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 4908 5556 4936 5596
rect 4985 5593 4997 5627
rect 5031 5624 5043 5627
rect 5644 5624 5672 5664
rect 5721 5661 5733 5695
rect 5767 5692 5779 5695
rect 5810 5692 5816 5704
rect 5767 5664 5816 5692
rect 5767 5661 5779 5664
rect 5721 5655 5779 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 5994 5652 6000 5704
rect 6052 5652 6058 5704
rect 6104 5701 6132 5732
rect 8220 5732 9220 5760
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 6380 5624 6408 5655
rect 7098 5652 7104 5704
rect 7156 5692 7162 5704
rect 7193 5695 7251 5701
rect 7193 5692 7205 5695
rect 7156 5664 7205 5692
rect 7156 5652 7162 5664
rect 7193 5661 7205 5664
rect 7239 5661 7251 5695
rect 7193 5655 7251 5661
rect 7282 5652 7288 5704
rect 7340 5652 7346 5704
rect 7374 5652 7380 5704
rect 7432 5692 7438 5704
rect 7469 5695 7527 5701
rect 7469 5692 7481 5695
rect 7432 5664 7481 5692
rect 7432 5652 7438 5664
rect 7469 5661 7481 5664
rect 7515 5661 7527 5695
rect 7469 5655 7527 5661
rect 5031 5596 5212 5624
rect 5644 5596 6408 5624
rect 7484 5624 7512 5655
rect 7558 5652 7564 5704
rect 7616 5652 7622 5704
rect 8220 5701 8248 5732
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 9766 5720 9772 5772
rect 9824 5760 9830 5772
rect 9824 5732 11100 5760
rect 9824 5720 9830 5732
rect 8205 5695 8263 5701
rect 8205 5661 8217 5695
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8570 5692 8576 5704
rect 8343 5664 8576 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10413 5695 10471 5701
rect 10413 5692 10425 5695
rect 10284 5664 10425 5692
rect 10284 5652 10290 5664
rect 10413 5661 10425 5664
rect 10459 5661 10471 5695
rect 10413 5655 10471 5661
rect 10502 5652 10508 5704
rect 10560 5652 10566 5704
rect 10689 5695 10747 5701
rect 10689 5661 10701 5695
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 8481 5627 8539 5633
rect 7484 5596 7880 5624
rect 5031 5593 5043 5596
rect 4985 5587 5043 5593
rect 5184 5568 5212 5596
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 4908 5528 5089 5556
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5077 5519 5135 5525
rect 5166 5516 5172 5568
rect 5224 5516 5230 5568
rect 5261 5559 5319 5565
rect 5261 5525 5273 5559
rect 5307 5556 5319 5559
rect 5626 5556 5632 5568
rect 5307 5528 5632 5556
rect 5307 5525 5319 5528
rect 5261 5519 5319 5525
rect 5626 5516 5632 5528
rect 5684 5556 5690 5568
rect 6270 5556 6276 5568
rect 5684 5528 6276 5556
rect 5684 5516 5690 5528
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 7742 5516 7748 5568
rect 7800 5516 7806 5568
rect 7852 5556 7880 5596
rect 8481 5593 8493 5627
rect 8527 5624 8539 5627
rect 8662 5624 8668 5636
rect 8527 5596 8668 5624
rect 8527 5593 8539 5596
rect 8481 5587 8539 5593
rect 8662 5584 8668 5596
rect 8720 5584 8726 5636
rect 10134 5584 10140 5636
rect 10192 5624 10198 5636
rect 10704 5624 10732 5655
rect 10778 5652 10784 5704
rect 10836 5652 10842 5704
rect 11072 5701 11100 5732
rect 11256 5701 11284 5800
rect 11330 5720 11336 5772
rect 11388 5760 11394 5772
rect 11885 5763 11943 5769
rect 11885 5760 11897 5763
rect 11388 5732 11897 5760
rect 11388 5720 11394 5732
rect 11885 5729 11897 5732
rect 11931 5729 11943 5763
rect 11885 5723 11943 5729
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 11241 5695 11299 5701
rect 11241 5661 11253 5695
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 12158 5652 12164 5704
rect 12216 5652 12222 5704
rect 10192 5596 10732 5624
rect 10192 5584 10198 5596
rect 10152 5556 10180 5584
rect 7852 5528 10180 5556
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 10965 5559 11023 5565
rect 10965 5556 10977 5559
rect 10744 5528 10977 5556
rect 10744 5516 10750 5528
rect 10965 5525 10977 5528
rect 11011 5525 11023 5559
rect 10965 5519 11023 5525
rect 1104 5466 12512 5488
rect 1104 5414 3036 5466
rect 3088 5414 3100 5466
rect 3152 5414 3164 5466
rect 3216 5414 3228 5466
rect 3280 5414 3292 5466
rect 3344 5414 5888 5466
rect 5940 5414 5952 5466
rect 6004 5414 6016 5466
rect 6068 5414 6080 5466
rect 6132 5414 6144 5466
rect 6196 5414 8740 5466
rect 8792 5414 8804 5466
rect 8856 5414 8868 5466
rect 8920 5414 8932 5466
rect 8984 5414 8996 5466
rect 9048 5414 11592 5466
rect 11644 5414 11656 5466
rect 11708 5414 11720 5466
rect 11772 5414 11784 5466
rect 11836 5414 11848 5466
rect 11900 5414 12512 5466
rect 1104 5392 12512 5414
rect 2593 5355 2651 5361
rect 2593 5321 2605 5355
rect 2639 5352 2651 5355
rect 4062 5352 4068 5364
rect 2639 5324 4068 5352
rect 2639 5321 2651 5324
rect 2593 5315 2651 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 7193 5355 7251 5361
rect 7193 5321 7205 5355
rect 7239 5352 7251 5355
rect 7282 5352 7288 5364
rect 7239 5324 7288 5352
rect 7239 5321 7251 5324
rect 7193 5315 7251 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 10502 5352 10508 5364
rect 8803 5324 10508 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 12066 5312 12072 5364
rect 12124 5312 12130 5364
rect 1673 5287 1731 5293
rect 1673 5253 1685 5287
rect 1719 5284 1731 5287
rect 2222 5284 2228 5296
rect 1719 5256 2228 5284
rect 1719 5253 1731 5256
rect 1673 5247 1731 5253
rect 2222 5244 2228 5256
rect 2280 5284 2286 5296
rect 4430 5284 4436 5296
rect 2280 5256 4436 5284
rect 2280 5244 2286 5256
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1489 5219 1547 5225
rect 1489 5216 1501 5219
rect 900 5188 1501 5216
rect 900 5176 906 5188
rect 1489 5185 1501 5188
rect 1535 5185 1547 5219
rect 1489 5179 1547 5185
rect 2501 5219 2559 5225
rect 2501 5185 2513 5219
rect 2547 5216 2559 5219
rect 2774 5216 2780 5228
rect 2547 5188 2780 5216
rect 2547 5185 2559 5188
rect 2501 5179 2559 5185
rect 2774 5176 2780 5188
rect 2832 5216 2838 5228
rect 3234 5216 3240 5228
rect 2832 5188 3240 5216
rect 2832 5176 2838 5188
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3510 5176 3516 5228
rect 3568 5176 3574 5228
rect 4080 5225 4108 5256
rect 4430 5244 4436 5256
rect 4488 5244 4494 5296
rect 5074 5244 5080 5296
rect 5132 5284 5138 5296
rect 5445 5287 5503 5293
rect 5445 5284 5457 5287
rect 5132 5256 5457 5284
rect 5132 5244 5138 5256
rect 5445 5253 5457 5256
rect 5491 5284 5503 5287
rect 8570 5284 8576 5296
rect 5491 5256 8576 5284
rect 5491 5253 5503 5256
rect 5445 5247 5503 5253
rect 8570 5244 8576 5256
rect 8628 5244 8634 5296
rect 11422 5244 11428 5296
rect 11480 5284 11486 5296
rect 11480 5256 11928 5284
rect 11480 5244 11486 5256
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4798 5176 4804 5228
rect 4856 5216 4862 5228
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 4856 5188 5273 5216
rect 4856 5176 4862 5188
rect 5261 5185 5273 5188
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 7469 5219 7527 5225
rect 7469 5216 7481 5219
rect 7156 5188 7481 5216
rect 7156 5176 7162 5188
rect 7469 5185 7481 5188
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 7926 5216 7932 5228
rect 7607 5188 7932 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 8389 5219 8447 5225
rect 8389 5185 8401 5219
rect 8435 5216 8447 5219
rect 9950 5216 9956 5228
rect 8435 5188 9956 5216
rect 8435 5185 8447 5188
rect 8389 5179 8447 5185
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 11900 5225 11928 5256
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 10192 5188 11529 5216
rect 10192 5176 10198 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 3881 5151 3939 5157
rect 3881 5148 3893 5151
rect 2096 5120 3893 5148
rect 2096 5108 2102 5120
rect 3881 5117 3893 5120
rect 3927 5148 3939 5151
rect 4249 5151 4307 5157
rect 4249 5148 4261 5151
rect 3927 5120 4261 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 4249 5117 4261 5120
rect 4295 5117 4307 5151
rect 4249 5111 4307 5117
rect 4525 5151 4583 5157
rect 4525 5117 4537 5151
rect 4571 5148 4583 5151
rect 6546 5148 6552 5160
rect 4571 5120 6552 5148
rect 4571 5117 4583 5120
rect 4525 5111 4583 5117
rect 6546 5108 6552 5120
rect 6604 5108 6610 5160
rect 7190 5108 7196 5160
rect 7248 5148 7254 5160
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 7248 5120 7389 5148
rect 7248 5108 7254 5120
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 7392 5080 7420 5111
rect 7650 5108 7656 5160
rect 7708 5108 7714 5160
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 8297 5151 8355 5157
rect 8297 5148 8309 5151
rect 7892 5120 8309 5148
rect 7892 5108 7898 5120
rect 8297 5117 8309 5120
rect 8343 5117 8355 5151
rect 8297 5111 8355 5117
rect 8478 5108 8484 5160
rect 8536 5108 8542 5160
rect 8573 5151 8631 5157
rect 8573 5117 8585 5151
rect 8619 5117 8631 5151
rect 8573 5111 8631 5117
rect 8588 5080 8616 5111
rect 7392 5052 8616 5080
rect 7006 4972 7012 5024
rect 7064 4972 7070 5024
rect 11698 4972 11704 5024
rect 11756 4972 11762 5024
rect 1104 4922 12512 4944
rect 1104 4870 2376 4922
rect 2428 4870 2440 4922
rect 2492 4870 2504 4922
rect 2556 4870 2568 4922
rect 2620 4870 2632 4922
rect 2684 4870 5228 4922
rect 5280 4870 5292 4922
rect 5344 4870 5356 4922
rect 5408 4870 5420 4922
rect 5472 4870 5484 4922
rect 5536 4870 8080 4922
rect 8132 4870 8144 4922
rect 8196 4870 8208 4922
rect 8260 4870 8272 4922
rect 8324 4870 8336 4922
rect 8388 4870 10932 4922
rect 10984 4870 10996 4922
rect 11048 4870 11060 4922
rect 11112 4870 11124 4922
rect 11176 4870 11188 4922
rect 11240 4870 12512 4922
rect 1104 4848 12512 4870
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2924 4780 2973 4808
rect 2924 4768 2930 4780
rect 2961 4777 2973 4780
rect 3007 4777 3019 4811
rect 2961 4771 3019 4777
rect 3234 4768 3240 4820
rect 3292 4808 3298 4820
rect 4062 4808 4068 4820
rect 3292 4780 4068 4808
rect 3292 4768 3298 4780
rect 4062 4768 4068 4780
rect 4120 4808 4126 4820
rect 4341 4811 4399 4817
rect 4341 4808 4353 4811
rect 4120 4780 4353 4808
rect 4120 4768 4126 4780
rect 4341 4777 4353 4780
rect 4387 4777 4399 4811
rect 4341 4771 4399 4777
rect 4798 4768 4804 4820
rect 4856 4768 4862 4820
rect 7193 4811 7251 4817
rect 7193 4777 7205 4811
rect 7239 4808 7251 4811
rect 7650 4808 7656 4820
rect 7239 4780 7656 4808
rect 7239 4777 7251 4780
rect 7193 4771 7251 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 7834 4768 7840 4820
rect 7892 4808 7898 4820
rect 8205 4811 8263 4817
rect 8205 4808 8217 4811
rect 7892 4780 8217 4808
rect 7892 4768 7898 4780
rect 8205 4777 8217 4780
rect 8251 4777 8263 4811
rect 8205 4771 8263 4777
rect 8478 4768 8484 4820
rect 8536 4808 8542 4820
rect 8536 4780 9076 4808
rect 8536 4768 8542 4780
rect 8113 4743 8171 4749
rect 8113 4740 8125 4743
rect 7576 4712 8125 4740
rect 4430 4632 4436 4684
rect 4488 4672 4494 4684
rect 4525 4675 4583 4681
rect 4525 4672 4537 4675
rect 4488 4644 4537 4672
rect 4488 4632 4494 4644
rect 4525 4641 4537 4644
rect 4571 4641 4583 4675
rect 4525 4635 4583 4641
rect 2222 4564 2228 4616
rect 2280 4604 2286 4616
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2280 4576 2881 4604
rect 2280 4564 2286 4576
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 3510 4604 3516 4616
rect 3099 4576 3516 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3510 4564 3516 4576
rect 3568 4604 3574 4616
rect 4154 4604 4160 4616
rect 3568 4576 4160 4604
rect 3568 4564 3574 4576
rect 4154 4564 4160 4576
rect 4212 4604 4218 4616
rect 4249 4607 4307 4613
rect 4249 4604 4261 4607
rect 4212 4576 4261 4604
rect 4212 4564 4218 4576
rect 4249 4573 4261 4576
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4982 4564 4988 4616
rect 5040 4564 5046 4616
rect 5074 4564 5080 4616
rect 5132 4604 5138 4616
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 5132 4576 5181 4604
rect 5132 4564 5138 4576
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 6362 4564 6368 4616
rect 6420 4604 6426 4616
rect 7377 4607 7435 4613
rect 7377 4604 7389 4607
rect 6420 4576 7389 4604
rect 6420 4564 6426 4576
rect 5077 4471 5135 4477
rect 5077 4437 5089 4471
rect 5123 4468 5135 4471
rect 5626 4468 5632 4480
rect 5123 4440 5632 4468
rect 5123 4437 5135 4440
rect 5077 4431 5135 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 7024 4468 7052 4576
rect 7377 4573 7389 4576
rect 7423 4573 7435 4607
rect 7377 4567 7435 4573
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4604 7527 4607
rect 7576 4604 7604 4712
rect 8113 4709 8125 4712
rect 8159 4709 8171 4743
rect 8941 4743 8999 4749
rect 8941 4740 8953 4743
rect 8113 4703 8171 4709
rect 8588 4712 8953 4740
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4672 7711 4675
rect 7699 4644 7880 4672
rect 7699 4641 7711 4644
rect 7653 4635 7711 4641
rect 7515 4576 7604 4604
rect 7515 4573 7527 4576
rect 7469 4567 7527 4573
rect 7098 4496 7104 4548
rect 7156 4536 7162 4548
rect 7668 4536 7696 4635
rect 7852 4613 7880 4644
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4573 7895 4607
rect 7837 4567 7895 4573
rect 7156 4508 7696 4536
rect 7760 4536 7788 4567
rect 7926 4564 7932 4616
rect 7984 4564 7990 4616
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8294 4604 8300 4616
rect 8159 4576 8300 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4604 8539 4607
rect 8588 4604 8616 4712
rect 8941 4709 8953 4712
rect 8987 4709 8999 4743
rect 8941 4703 8999 4709
rect 8665 4675 8723 4681
rect 8665 4641 8677 4675
rect 8711 4672 8723 4675
rect 9048 4672 9076 4780
rect 10134 4768 10140 4820
rect 10192 4768 10198 4820
rect 10686 4768 10692 4820
rect 10744 4768 10750 4820
rect 10965 4811 11023 4817
rect 10965 4777 10977 4811
rect 11011 4808 11023 4811
rect 11974 4808 11980 4820
rect 11011 4780 11980 4808
rect 11011 4777 11023 4780
rect 10965 4771 11023 4777
rect 10318 4700 10324 4752
rect 10376 4740 10382 4752
rect 10980 4740 11008 4771
rect 11974 4768 11980 4780
rect 12032 4768 12038 4820
rect 10376 4712 11008 4740
rect 10376 4700 10382 4712
rect 8711 4644 9260 4672
rect 8711 4641 8723 4644
rect 8665 4635 8723 4641
rect 9232 4613 9260 4644
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 10468 4644 10916 4672
rect 10468 4632 10474 4644
rect 8527 4576 8616 4604
rect 8757 4607 8815 4613
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 8757 4573 8769 4607
rect 8803 4604 8815 4607
rect 9217 4607 9275 4613
rect 8803 4576 9168 4604
rect 8803 4573 8815 4576
rect 8757 4567 8815 4573
rect 7944 4536 7972 4564
rect 7760 4508 7972 4536
rect 7156 4496 7162 4508
rect 8404 4468 8432 4567
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 9140 4545 9168 4576
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9398 4604 9404 4616
rect 9263 4576 9404 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 9950 4564 9956 4616
rect 10008 4604 10014 4616
rect 10888 4613 10916 4644
rect 10962 4632 10968 4684
rect 11020 4672 11026 4684
rect 11149 4675 11207 4681
rect 11149 4672 11161 4675
rect 11020 4644 11161 4672
rect 11020 4632 11026 4644
rect 11149 4641 11161 4644
rect 11195 4641 11207 4675
rect 11149 4635 11207 4641
rect 10262 4607 10320 4613
rect 10262 4604 10274 4607
rect 10008 4576 10274 4604
rect 10008 4564 10014 4576
rect 10262 4573 10274 4576
rect 10308 4573 10320 4607
rect 10262 4567 10320 4573
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 8941 4539 8999 4545
rect 8941 4536 8953 4539
rect 8628 4508 8953 4536
rect 8628 4496 8634 4508
rect 8941 4505 8953 4508
rect 8987 4505 8999 4539
rect 8941 4499 8999 4505
rect 9125 4539 9183 4545
rect 9125 4505 9137 4539
rect 9171 4536 9183 4539
rect 9968 4536 9996 4564
rect 9171 4508 9996 4536
rect 10796 4536 10824 4567
rect 11514 4536 11520 4548
rect 10796 4508 11520 4536
rect 9171 4505 9183 4508
rect 9125 4499 9183 4505
rect 11514 4496 11520 4508
rect 11572 4496 11578 4548
rect 7024 4440 8432 4468
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10321 4471 10379 4477
rect 10321 4468 10333 4471
rect 10284 4440 10333 4468
rect 10284 4428 10290 4440
rect 10321 4437 10333 4440
rect 10367 4437 10379 4471
rect 10321 4431 10379 4437
rect 11146 4428 11152 4480
rect 11204 4428 11210 4480
rect 1104 4378 12512 4400
rect 1104 4326 3036 4378
rect 3088 4326 3100 4378
rect 3152 4326 3164 4378
rect 3216 4326 3228 4378
rect 3280 4326 3292 4378
rect 3344 4326 5888 4378
rect 5940 4326 5952 4378
rect 6004 4326 6016 4378
rect 6068 4326 6080 4378
rect 6132 4326 6144 4378
rect 6196 4326 8740 4378
rect 8792 4326 8804 4378
rect 8856 4326 8868 4378
rect 8920 4326 8932 4378
rect 8984 4326 8996 4378
rect 9048 4326 11592 4378
rect 11644 4326 11656 4378
rect 11708 4326 11720 4378
rect 11772 4326 11784 4378
rect 11836 4326 11848 4378
rect 11900 4326 12512 4378
rect 1104 4304 12512 4326
rect 4430 4264 4436 4276
rect 3896 4236 4436 4264
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4128 3847 4131
rect 3896 4128 3924 4236
rect 4430 4224 4436 4236
rect 4488 4224 4494 4276
rect 5534 4264 5540 4276
rect 5460 4236 5540 4264
rect 4062 4156 4068 4208
rect 4120 4196 4126 4208
rect 4157 4199 4215 4205
rect 4157 4196 4169 4199
rect 4120 4168 4169 4196
rect 4120 4156 4126 4168
rect 4157 4165 4169 4168
rect 4203 4165 4215 4199
rect 4157 4159 4215 4165
rect 4982 4156 4988 4208
rect 5040 4156 5046 4208
rect 3835 4100 3924 4128
rect 3835 4097 3847 4100
rect 3789 4091 3847 4097
rect 4338 4088 4344 4140
rect 4396 4128 4402 4140
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4396 4100 4905 4128
rect 4396 4088 4402 4100
rect 4893 4097 4905 4100
rect 4939 4097 4951 4131
rect 5000 4128 5028 4156
rect 5353 4131 5411 4137
rect 5353 4128 5365 4131
rect 5000 4100 5365 4128
rect 4893 4091 4951 4097
rect 5353 4097 5365 4100
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 4430 4020 4436 4072
rect 4488 4060 4494 4072
rect 4709 4063 4767 4069
rect 4709 4060 4721 4063
rect 4488 4032 4721 4060
rect 4488 4020 4494 4032
rect 4709 4029 4721 4032
rect 4755 4029 4767 4063
rect 4709 4023 4767 4029
rect 4798 4020 4804 4072
rect 4856 4020 4862 4072
rect 4154 3884 4160 3936
rect 4212 3884 4218 3936
rect 4338 3884 4344 3936
rect 4396 3884 4402 3936
rect 4525 3927 4583 3933
rect 4525 3893 4537 3927
rect 4571 3924 4583 3927
rect 4614 3924 4620 3936
rect 4571 3896 4620 3924
rect 4571 3893 4583 3896
rect 4525 3887 4583 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4908 3924 4936 4091
rect 4985 4063 5043 4069
rect 4985 4029 4997 4063
rect 5031 4029 5043 4063
rect 4985 4023 5043 4029
rect 5000 3992 5028 4023
rect 5074 4020 5080 4072
rect 5132 4060 5138 4072
rect 5261 4063 5319 4069
rect 5261 4060 5273 4063
rect 5132 4032 5273 4060
rect 5132 4020 5138 4032
rect 5261 4029 5273 4032
rect 5307 4029 5319 4063
rect 5261 4023 5319 4029
rect 5460 3992 5488 4236
rect 5534 4224 5540 4236
rect 5592 4264 5598 4276
rect 8021 4267 8079 4273
rect 8021 4264 8033 4267
rect 5592 4236 8033 4264
rect 5592 4224 5598 4236
rect 8021 4233 8033 4236
rect 8067 4264 8079 4267
rect 10226 4264 10232 4276
rect 8067 4236 10232 4264
rect 8067 4233 8079 4236
rect 8021 4227 8079 4233
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 5718 4156 5724 4208
rect 5776 4196 5782 4208
rect 5965 4199 6023 4205
rect 5965 4196 5977 4199
rect 5776 4168 5977 4196
rect 5776 4156 5782 4168
rect 5965 4165 5977 4168
rect 6011 4165 6023 4199
rect 5965 4159 6023 4165
rect 6181 4199 6239 4205
rect 6181 4165 6193 4199
rect 6227 4165 6239 4199
rect 6181 4159 6239 4165
rect 9677 4199 9735 4205
rect 9677 4165 9689 4199
rect 9723 4196 9735 4199
rect 10134 4196 10140 4208
rect 9723 4168 10140 4196
rect 9723 4165 9735 4168
rect 9677 4159 9735 4165
rect 6196 4128 6224 4159
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 10410 4196 10416 4208
rect 10244 4168 10416 4196
rect 6822 4128 6828 4140
rect 5000 3964 5488 3992
rect 5644 4100 6828 4128
rect 5644 3924 5672 4100
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 7742 4128 7748 4140
rect 7699 4100 7748 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 10244 4137 10272 4168
rect 10410 4156 10416 4168
rect 10468 4196 10474 4208
rect 10686 4196 10692 4208
rect 10468 4168 10692 4196
rect 10468 4156 10474 4168
rect 10686 4156 10692 4168
rect 10744 4196 10750 4208
rect 10744 4168 10916 4196
rect 10744 4156 10750 4168
rect 8024 4131 8082 4137
rect 8024 4128 8036 4131
rect 7984 4100 8036 4128
rect 7984 4088 7990 4100
rect 8024 4097 8036 4100
rect 8070 4097 8082 4131
rect 8024 4091 8082 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4128 9919 4131
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9907 4100 10057 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 10318 4088 10324 4140
rect 10376 4088 10382 4140
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 5721 4063 5779 4069
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 6362 4060 6368 4072
rect 5767 4032 6368 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 6362 4020 6368 4032
rect 6420 4020 6426 4072
rect 7558 4020 7564 4072
rect 7616 4020 7622 4072
rect 10520 4060 10548 4091
rect 10594 4088 10600 4140
rect 10652 4128 10658 4140
rect 10781 4131 10839 4137
rect 10781 4128 10793 4131
rect 10652 4100 10793 4128
rect 10652 4088 10658 4100
rect 10781 4097 10793 4100
rect 10827 4097 10839 4131
rect 10888 4128 10916 4168
rect 11146 4156 11152 4208
rect 11204 4196 11210 4208
rect 11204 4168 11836 4196
rect 11204 4156 11210 4168
rect 11808 4137 11836 4168
rect 11057 4131 11115 4137
rect 11057 4128 11069 4131
rect 10888 4100 11069 4128
rect 10781 4091 10839 4097
rect 11057 4097 11069 4100
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 11241 4131 11299 4137
rect 11241 4097 11253 4131
rect 11287 4128 11299 4131
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11287 4100 11713 4128
rect 11287 4097 11299 4100
rect 11241 4091 11299 4097
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 10060 4032 10548 4060
rect 10060 4004 10088 4032
rect 11514 4020 11520 4072
rect 11572 4020 11578 4072
rect 5810 3952 5816 4004
rect 5868 3952 5874 4004
rect 10042 3952 10048 4004
rect 10100 3952 10106 4004
rect 10410 3952 10416 4004
rect 10468 3952 10474 4004
rect 10778 3952 10784 4004
rect 10836 3992 10842 4004
rect 10873 3995 10931 4001
rect 10873 3992 10885 3995
rect 10836 3964 10885 3992
rect 10836 3952 10842 3964
rect 10873 3961 10885 3964
rect 10919 3961 10931 3995
rect 10873 3955 10931 3961
rect 10965 3995 11023 4001
rect 10965 3961 10977 3995
rect 11011 3961 11023 3995
rect 10965 3955 11023 3961
rect 4908 3896 5672 3924
rect 5994 3884 6000 3936
rect 6052 3884 6058 3936
rect 8205 3927 8263 3933
rect 8205 3893 8217 3927
rect 8251 3924 8263 3927
rect 8478 3924 8484 3936
rect 8251 3896 8484 3924
rect 8251 3893 8263 3896
rect 8205 3887 8263 3893
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9493 3927 9551 3933
rect 9493 3924 9505 3927
rect 9272 3896 9505 3924
rect 9272 3884 9278 3896
rect 9493 3893 9505 3896
rect 9539 3893 9551 3927
rect 9493 3887 9551 3893
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 10980 3924 11008 3955
rect 10376 3896 11008 3924
rect 10376 3884 10382 3896
rect 1104 3834 12512 3856
rect 1104 3782 2376 3834
rect 2428 3782 2440 3834
rect 2492 3782 2504 3834
rect 2556 3782 2568 3834
rect 2620 3782 2632 3834
rect 2684 3782 5228 3834
rect 5280 3782 5292 3834
rect 5344 3782 5356 3834
rect 5408 3782 5420 3834
rect 5472 3782 5484 3834
rect 5536 3782 8080 3834
rect 8132 3782 8144 3834
rect 8196 3782 8208 3834
rect 8260 3782 8272 3834
rect 8324 3782 8336 3834
rect 8388 3782 10932 3834
rect 10984 3782 10996 3834
rect 11048 3782 11060 3834
rect 11112 3782 11124 3834
rect 11176 3782 11188 3834
rect 11240 3782 12512 3834
rect 1104 3760 12512 3782
rect 4430 3680 4436 3732
rect 4488 3680 4494 3732
rect 4709 3723 4767 3729
rect 4709 3689 4721 3723
rect 4755 3689 4767 3723
rect 4709 3683 4767 3689
rect 4341 3655 4399 3661
rect 4341 3621 4353 3655
rect 4387 3652 4399 3655
rect 4724 3652 4752 3683
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 5261 3723 5319 3729
rect 5261 3720 5273 3723
rect 4856 3692 5273 3720
rect 4856 3680 4862 3692
rect 5261 3689 5273 3692
rect 5307 3689 5319 3723
rect 5261 3683 5319 3689
rect 5994 3680 6000 3732
rect 6052 3680 6058 3732
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 10410 3720 10416 3732
rect 9723 3692 10416 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 10410 3680 10416 3692
rect 10468 3680 10474 3732
rect 4387 3624 5580 3652
rect 4387 3621 4399 3624
rect 4341 3615 4399 3621
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 4632 3556 5457 3584
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4338 3476 4344 3528
rect 4396 3476 4402 3528
rect 4430 3476 4436 3528
rect 4488 3516 4494 3528
rect 4632 3525 4660 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 4488 3488 4629 3516
rect 4488 3476 4494 3488
rect 4617 3485 4629 3488
rect 4663 3485 4675 3519
rect 4985 3519 5043 3525
rect 4985 3515 4997 3519
rect 4617 3479 4675 3485
rect 4908 3487 4997 3515
rect 4908 3448 4936 3487
rect 4985 3485 4997 3487
rect 5031 3485 5043 3519
rect 4985 3479 5043 3485
rect 5077 3519 5135 3525
rect 5077 3485 5089 3519
rect 5123 3515 5135 3519
rect 5350 3516 5356 3528
rect 5181 3515 5356 3516
rect 5123 3488 5356 3515
rect 5123 3487 5209 3488
rect 5123 3485 5135 3487
rect 5077 3479 5135 3485
rect 5350 3476 5356 3488
rect 5408 3476 5414 3528
rect 5552 3525 5580 3624
rect 5626 3612 5632 3664
rect 5684 3652 5690 3664
rect 6454 3652 6460 3664
rect 5684 3624 5948 3652
rect 5684 3612 5690 3624
rect 5718 3544 5724 3596
rect 5776 3584 5782 3596
rect 5920 3593 5948 3624
rect 6104 3624 6460 3652
rect 5813 3587 5871 3593
rect 5813 3584 5825 3587
rect 5776 3556 5825 3584
rect 5776 3544 5782 3556
rect 5813 3553 5825 3556
rect 5859 3553 5871 3587
rect 5813 3547 5871 3553
rect 5905 3587 5963 3593
rect 5905 3553 5917 3587
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 6104 3525 6132 3624
rect 6454 3612 6460 3624
rect 6512 3652 6518 3664
rect 9306 3652 9312 3664
rect 6512 3624 9312 3652
rect 6512 3612 6518 3624
rect 9306 3612 9312 3624
rect 9364 3612 9370 3664
rect 9585 3655 9643 3661
rect 9585 3621 9597 3655
rect 9631 3652 9643 3655
rect 9950 3652 9956 3664
rect 9631 3624 9956 3652
rect 9631 3621 9643 3624
rect 9585 3615 9643 3621
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 6733 3587 6791 3593
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 6914 3584 6920 3596
rect 6779 3556 6920 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 6914 3544 6920 3556
rect 6972 3584 6978 3596
rect 7285 3587 7343 3593
rect 7285 3584 7297 3587
rect 6972 3556 7297 3584
rect 6972 3544 6978 3556
rect 7285 3553 7297 3556
rect 7331 3553 7343 3587
rect 8021 3587 8079 3593
rect 8021 3584 8033 3587
rect 7285 3547 7343 3553
rect 7484 3556 8033 3584
rect 7484 3528 7512 3556
rect 8021 3553 8033 3556
rect 8067 3553 8079 3587
rect 8021 3547 8079 3553
rect 8481 3587 8539 3593
rect 8481 3553 8493 3587
rect 8527 3584 8539 3587
rect 9217 3587 9275 3593
rect 9217 3584 9229 3587
rect 8527 3556 9229 3584
rect 8527 3553 8539 3556
rect 8481 3547 8539 3553
rect 9217 3553 9229 3556
rect 9263 3584 9275 3587
rect 9766 3584 9772 3596
rect 9263 3556 9772 3584
rect 9263 3553 9275 3556
rect 9217 3547 9275 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 10428 3584 10456 3680
rect 10428 3556 11008 3584
rect 5537 3519 5595 3525
rect 5537 3485 5549 3519
rect 5583 3485 5595 3519
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 5537 3479 5595 3485
rect 5828 3488 6009 3516
rect 5828 3460 5856 3488
rect 5997 3485 6009 3488
rect 6043 3485 6055 3519
rect 5997 3479 6055 3485
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3485 6147 3519
rect 6089 3479 6147 3485
rect 6549 3519 6607 3525
rect 6549 3485 6561 3519
rect 6595 3485 6607 3519
rect 6549 3479 6607 3485
rect 6825 3519 6883 3525
rect 6825 3485 6837 3519
rect 6871 3516 6883 3519
rect 7098 3516 7104 3528
rect 6871 3488 7104 3516
rect 6871 3485 6883 3488
rect 6825 3479 6883 3485
rect 5718 3448 5724 3460
rect 4908 3420 5724 3448
rect 5718 3408 5724 3420
rect 5776 3408 5782 3460
rect 5810 3408 5816 3460
rect 5868 3408 5874 3460
rect 6270 3408 6276 3460
rect 6328 3408 6334 3460
rect 6564 3448 6592 3479
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7466 3476 7472 3528
rect 7524 3476 7530 3528
rect 7745 3519 7803 3525
rect 7745 3485 7757 3519
rect 7791 3485 7803 3519
rect 7745 3479 7803 3485
rect 8113 3519 8171 3525
rect 8113 3485 8125 3519
rect 8159 3516 8171 3519
rect 9398 3516 9404 3528
rect 8159 3488 9404 3516
rect 8159 3485 8171 3488
rect 8113 3479 8171 3485
rect 7006 3448 7012 3460
rect 6564 3420 7012 3448
rect 7006 3408 7012 3420
rect 7064 3448 7070 3460
rect 7760 3448 7788 3479
rect 7064 3420 7788 3448
rect 7064 3408 7070 3420
rect 6365 3383 6423 3389
rect 6365 3349 6377 3383
rect 6411 3380 6423 3383
rect 6546 3380 6552 3392
rect 6411 3352 6552 3380
rect 6411 3349 6423 3352
rect 6365 3343 6423 3349
rect 6546 3340 6552 3352
rect 6604 3340 6610 3392
rect 7653 3383 7711 3389
rect 7653 3349 7665 3383
rect 7699 3380 7711 3383
rect 8128 3380 8156 3479
rect 9398 3476 9404 3488
rect 9456 3476 9462 3528
rect 10042 3476 10048 3528
rect 10100 3476 10106 3528
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 10318 3476 10324 3528
rect 10376 3516 10382 3528
rect 10980 3525 11008 3556
rect 10505 3519 10563 3525
rect 10505 3516 10517 3519
rect 10376 3488 10517 3516
rect 10376 3476 10382 3488
rect 10505 3485 10517 3488
rect 10551 3485 10563 3519
rect 10505 3479 10563 3485
rect 10965 3519 11023 3525
rect 10965 3485 10977 3519
rect 11011 3485 11023 3519
rect 10965 3479 11023 3485
rect 11333 3519 11391 3525
rect 11333 3485 11345 3519
rect 11379 3485 11391 3519
rect 11333 3479 11391 3485
rect 9306 3408 9312 3460
rect 9364 3448 9370 3460
rect 9769 3451 9827 3457
rect 9769 3448 9781 3451
rect 9364 3420 9781 3448
rect 9364 3408 9370 3420
rect 9769 3417 9781 3420
rect 9815 3417 9827 3451
rect 9769 3411 9827 3417
rect 10686 3408 10692 3460
rect 10744 3448 10750 3460
rect 11348 3448 11376 3479
rect 10744 3420 11376 3448
rect 10744 3408 10750 3420
rect 7699 3352 8156 3380
rect 7699 3349 7711 3352
rect 7653 3343 7711 3349
rect 1104 3290 12512 3312
rect 1104 3238 3036 3290
rect 3088 3238 3100 3290
rect 3152 3238 3164 3290
rect 3216 3238 3228 3290
rect 3280 3238 3292 3290
rect 3344 3238 5888 3290
rect 5940 3238 5952 3290
rect 6004 3238 6016 3290
rect 6068 3238 6080 3290
rect 6132 3238 6144 3290
rect 6196 3238 8740 3290
rect 8792 3238 8804 3290
rect 8856 3238 8868 3290
rect 8920 3238 8932 3290
rect 8984 3238 8996 3290
rect 9048 3238 11592 3290
rect 11644 3238 11656 3290
rect 11708 3238 11720 3290
rect 11772 3238 11784 3290
rect 11836 3238 11848 3290
rect 11900 3238 12512 3290
rect 1104 3216 12512 3238
rect 5074 3136 5080 3188
rect 5132 3176 5138 3188
rect 5261 3179 5319 3185
rect 5261 3176 5273 3179
rect 5132 3148 5273 3176
rect 5132 3136 5138 3148
rect 5261 3145 5273 3148
rect 5307 3145 5319 3179
rect 5261 3139 5319 3145
rect 5537 3179 5595 3185
rect 5537 3145 5549 3179
rect 5583 3176 5595 3179
rect 5718 3176 5724 3188
rect 5583 3148 5724 3176
rect 5583 3145 5595 3148
rect 5537 3139 5595 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 5905 3179 5963 3185
rect 5905 3176 5917 3179
rect 5868 3148 5917 3176
rect 5868 3136 5874 3148
rect 5905 3145 5917 3148
rect 5951 3176 5963 3179
rect 7377 3179 7435 3185
rect 5951 3148 6316 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 6288 3108 6316 3148
rect 7377 3145 7389 3179
rect 7423 3145 7435 3179
rect 7377 3139 7435 3145
rect 7392 3108 7420 3139
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 9033 3179 9091 3185
rect 9033 3176 9045 3179
rect 7616 3148 9045 3176
rect 7616 3136 7622 3148
rect 9033 3145 9045 3148
rect 9079 3145 9091 3179
rect 9033 3139 9091 3145
rect 9201 3179 9259 3185
rect 9201 3145 9213 3179
rect 9247 3176 9259 3179
rect 9306 3176 9312 3188
rect 9247 3148 9312 3176
rect 9247 3145 9259 3148
rect 9201 3139 9259 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10229 3179 10287 3185
rect 10229 3176 10241 3179
rect 10100 3148 10241 3176
rect 10100 3136 10106 3148
rect 10229 3145 10241 3148
rect 10275 3145 10287 3179
rect 10229 3139 10287 3145
rect 7745 3111 7803 3117
rect 7745 3108 7757 3111
rect 5736 3080 6132 3108
rect 6288 3080 7144 3108
rect 7392 3080 7757 3108
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4706 3040 4712 3052
rect 4212 3012 4712 3040
rect 4212 3000 4218 3012
rect 4706 3000 4712 3012
rect 4764 3040 4770 3052
rect 4893 3043 4951 3049
rect 4893 3040 4905 3043
rect 4764 3012 4905 3040
rect 4764 3000 4770 3012
rect 4893 3009 4905 3012
rect 4939 3040 4951 3043
rect 5626 3040 5632 3052
rect 4939 3012 5632 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 5736 3049 5764 3080
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 5997 3043 6055 3049
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 6104 3040 6132 3080
rect 6270 3040 6276 3052
rect 6104 3012 6276 3040
rect 5997 3003 6055 3009
rect 4338 2932 4344 2984
rect 4396 2972 4402 2984
rect 4985 2975 5043 2981
rect 4985 2972 4997 2975
rect 4396 2944 4997 2972
rect 4396 2932 4402 2944
rect 4985 2941 4997 2944
rect 5031 2941 5043 2975
rect 6012 2972 6040 3003
rect 6270 3000 6276 3012
rect 6328 3000 6334 3052
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 7006 3000 7012 3052
rect 7064 3000 7070 3052
rect 6454 2972 6460 2984
rect 6012 2944 6460 2972
rect 4985 2935 5043 2941
rect 5000 2904 5028 2935
rect 6454 2932 6460 2944
rect 6512 2932 6518 2984
rect 6914 2932 6920 2984
rect 6972 2932 6978 2984
rect 7116 2972 7144 3080
rect 7484 3049 7512 3080
rect 7745 3077 7757 3080
rect 7791 3077 7803 3111
rect 9401 3111 9459 3117
rect 9401 3108 9413 3111
rect 7745 3071 7803 3077
rect 8404 3080 9413 3108
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7926 3040 7932 3052
rect 7699 3012 7932 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 8297 3043 8355 3049
rect 8297 3040 8309 3043
rect 8159 3012 8309 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 8297 3009 8309 3012
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7116 2944 7573 2972
rect 7561 2941 7573 2944
rect 7607 2972 7619 2975
rect 8205 2975 8263 2981
rect 8205 2972 8217 2975
rect 7607 2944 8217 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 8205 2941 8217 2944
rect 8251 2941 8263 2975
rect 8205 2935 8263 2941
rect 6546 2904 6552 2916
rect 5000 2876 6552 2904
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 6822 2864 6828 2916
rect 6880 2904 6886 2916
rect 8404 2904 8432 3080
rect 9401 3077 9413 3080
rect 9447 3108 9459 3111
rect 9858 3108 9864 3120
rect 9447 3080 9864 3108
rect 9447 3077 9459 3080
rect 9401 3071 9459 3077
rect 9858 3068 9864 3080
rect 9916 3108 9922 3120
rect 10244 3108 10272 3139
rect 10778 3136 10784 3188
rect 10836 3136 10842 3188
rect 9916 3080 10180 3108
rect 10244 3080 11008 3108
rect 9916 3068 9922 3080
rect 9766 3000 9772 3052
rect 9824 3000 9830 3052
rect 10152 3040 10180 3080
rect 10152 3012 10364 3040
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 10134 2972 10140 2984
rect 8803 2944 10140 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 10336 2972 10364 3012
rect 10410 3000 10416 3052
rect 10468 3040 10474 3052
rect 10980 3049 11008 3080
rect 10689 3043 10747 3049
rect 10689 3040 10701 3043
rect 10468 3012 10701 3040
rect 10468 3000 10474 3012
rect 10689 3009 10701 3012
rect 10735 3009 10747 3043
rect 10689 3003 10747 3009
rect 10873 3043 10931 3049
rect 10873 3009 10885 3043
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 10594 2972 10600 2984
rect 10336 2944 10600 2972
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10888 2972 10916 3003
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 10888 2944 11069 2972
rect 11057 2941 11069 2944
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 6880 2876 8432 2904
rect 6880 2864 6886 2876
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 6457 2839 6515 2845
rect 6457 2836 6469 2839
rect 6328 2808 6469 2836
rect 6328 2796 6334 2808
rect 6457 2805 6469 2808
rect 6503 2805 6515 2839
rect 6457 2799 6515 2805
rect 9214 2796 9220 2848
rect 9272 2796 9278 2848
rect 10042 2796 10048 2848
rect 10100 2796 10106 2848
rect 1104 2746 12512 2768
rect 1104 2694 2376 2746
rect 2428 2694 2440 2746
rect 2492 2694 2504 2746
rect 2556 2694 2568 2746
rect 2620 2694 2632 2746
rect 2684 2694 5228 2746
rect 5280 2694 5292 2746
rect 5344 2694 5356 2746
rect 5408 2694 5420 2746
rect 5472 2694 5484 2746
rect 5536 2694 8080 2746
rect 8132 2694 8144 2746
rect 8196 2694 8208 2746
rect 8260 2694 8272 2746
rect 8324 2694 8336 2746
rect 8388 2694 10932 2746
rect 10984 2694 10996 2746
rect 11048 2694 11060 2746
rect 11112 2694 11124 2746
rect 11176 2694 11188 2746
rect 11240 2694 12512 2746
rect 1104 2672 12512 2694
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 5040 2604 6653 2632
rect 5040 2592 5046 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 6641 2595 6699 2601
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 7984 2604 8493 2632
rect 7984 2592 7990 2604
rect 8481 2601 8493 2604
rect 8527 2601 8539 2635
rect 8481 2595 8539 2601
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10229 2635 10287 2641
rect 10229 2632 10241 2635
rect 10100 2604 10241 2632
rect 10100 2592 10106 2604
rect 10229 2601 10241 2604
rect 10275 2601 10287 2635
rect 10229 2595 10287 2601
rect 4341 2567 4399 2573
rect 4341 2533 4353 2567
rect 4387 2564 4399 2567
rect 5166 2564 5172 2576
rect 4387 2536 5172 2564
rect 4387 2533 4399 2536
rect 4341 2527 4399 2533
rect 5166 2524 5172 2536
rect 5224 2524 5230 2576
rect 5718 2456 5724 2508
rect 5776 2496 5782 2508
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5776 2468 5917 2496
rect 5776 2456 5782 2468
rect 5905 2465 5917 2468
rect 5951 2465 5963 2499
rect 5905 2459 5963 2465
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7469 2499 7527 2505
rect 7469 2496 7481 2499
rect 7064 2468 7481 2496
rect 7064 2456 7070 2468
rect 7469 2465 7481 2468
rect 7515 2465 7527 2499
rect 7469 2459 7527 2465
rect 9398 2456 9404 2508
rect 9456 2456 9462 2508
rect 4522 2388 4528 2440
rect 4580 2388 4586 2440
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6181 2431 6239 2437
rect 6181 2428 6193 2431
rect 5868 2400 6193 2428
rect 5868 2388 5874 2400
rect 6181 2397 6193 2400
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 7156 2400 7205 2428
rect 7156 2388 7162 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8478 2428 8484 2440
rect 8435 2400 8484 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 4893 2363 4951 2369
rect 4893 2360 4905 2363
rect 4540 2332 4905 2360
rect 4540 2304 4568 2332
rect 4893 2329 4905 2332
rect 4939 2329 4951 2363
rect 4893 2323 4951 2329
rect 6454 2320 6460 2372
rect 6512 2360 6518 2372
rect 6733 2363 6791 2369
rect 6733 2360 6745 2363
rect 6512 2332 6745 2360
rect 6512 2320 6518 2332
rect 6733 2329 6745 2332
rect 6779 2329 6791 2363
rect 8680 2360 8708 2391
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 10045 2431 10103 2437
rect 10045 2428 10057 2431
rect 9732 2400 10057 2428
rect 9732 2388 9738 2400
rect 10045 2397 10057 2400
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 6733 2323 6791 2329
rect 8404 2332 8708 2360
rect 8404 2304 8432 2332
rect 4522 2252 4528 2304
rect 4580 2252 4586 2304
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 8205 2295 8263 2301
rect 8205 2292 8217 2295
rect 7800 2264 8217 2292
rect 7800 2252 7806 2264
rect 8205 2261 8217 2264
rect 8251 2261 8263 2295
rect 8205 2255 8263 2261
rect 8386 2252 8392 2304
rect 8444 2252 8450 2304
rect 1104 2202 12512 2224
rect 1104 2150 3036 2202
rect 3088 2150 3100 2202
rect 3152 2150 3164 2202
rect 3216 2150 3228 2202
rect 3280 2150 3292 2202
rect 3344 2150 5888 2202
rect 5940 2150 5952 2202
rect 6004 2150 6016 2202
rect 6068 2150 6080 2202
rect 6132 2150 6144 2202
rect 6196 2150 8740 2202
rect 8792 2150 8804 2202
rect 8856 2150 8868 2202
rect 8920 2150 8932 2202
rect 8984 2150 8996 2202
rect 9048 2150 11592 2202
rect 11644 2150 11656 2202
rect 11708 2150 11720 2202
rect 11772 2150 11784 2202
rect 11836 2150 11848 2202
rect 11900 2150 12512 2202
rect 1104 2128 12512 2150
<< via1 >>
rect 2376 13574 2428 13626
rect 2440 13574 2492 13626
rect 2504 13574 2556 13626
rect 2568 13574 2620 13626
rect 2632 13574 2684 13626
rect 5228 13574 5280 13626
rect 5292 13574 5344 13626
rect 5356 13574 5408 13626
rect 5420 13574 5472 13626
rect 5484 13574 5536 13626
rect 8080 13574 8132 13626
rect 8144 13574 8196 13626
rect 8208 13574 8260 13626
rect 8272 13574 8324 13626
rect 8336 13574 8388 13626
rect 10932 13574 10984 13626
rect 10996 13574 11048 13626
rect 11060 13574 11112 13626
rect 11124 13574 11176 13626
rect 11188 13574 11240 13626
rect 7748 13336 7800 13388
rect 4528 13268 4580 13320
rect 6460 13268 6512 13320
rect 7104 13268 7156 13320
rect 7840 13200 7892 13252
rect 4620 13132 4672 13184
rect 6276 13132 6328 13184
rect 7196 13132 7248 13184
rect 3036 13030 3088 13082
rect 3100 13030 3152 13082
rect 3164 13030 3216 13082
rect 3228 13030 3280 13082
rect 3292 13030 3344 13082
rect 5888 13030 5940 13082
rect 5952 13030 6004 13082
rect 6016 13030 6068 13082
rect 6080 13030 6132 13082
rect 6144 13030 6196 13082
rect 8740 13030 8792 13082
rect 8804 13030 8856 13082
rect 8868 13030 8920 13082
rect 8932 13030 8984 13082
rect 8996 13030 9048 13082
rect 11592 13030 11644 13082
rect 11656 13030 11708 13082
rect 11720 13030 11772 13082
rect 11784 13030 11836 13082
rect 11848 13030 11900 13082
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 4988 12792 5040 12844
rect 7104 12792 7156 12844
rect 7656 12792 7708 12844
rect 9036 12835 9088 12844
rect 9036 12801 9045 12835
rect 9045 12801 9079 12835
rect 9079 12801 9088 12835
rect 9036 12792 9088 12801
rect 4804 12767 4856 12776
rect 4804 12733 4813 12767
rect 4813 12733 4847 12767
rect 4847 12733 4856 12767
rect 4804 12724 4856 12733
rect 5816 12724 5868 12776
rect 7932 12767 7984 12776
rect 7932 12733 7941 12767
rect 7941 12733 7975 12767
rect 7975 12733 7984 12767
rect 7932 12724 7984 12733
rect 8944 12724 8996 12776
rect 10324 12656 10376 12708
rect 1676 12588 1728 12640
rect 6736 12588 6788 12640
rect 10232 12588 10284 12640
rect 2376 12486 2428 12538
rect 2440 12486 2492 12538
rect 2504 12486 2556 12538
rect 2568 12486 2620 12538
rect 2632 12486 2684 12538
rect 5228 12486 5280 12538
rect 5292 12486 5344 12538
rect 5356 12486 5408 12538
rect 5420 12486 5472 12538
rect 5484 12486 5536 12538
rect 8080 12486 8132 12538
rect 8144 12486 8196 12538
rect 8208 12486 8260 12538
rect 8272 12486 8324 12538
rect 8336 12486 8388 12538
rect 10932 12486 10984 12538
rect 10996 12486 11048 12538
rect 11060 12486 11112 12538
rect 11124 12486 11176 12538
rect 11188 12486 11240 12538
rect 4712 12427 4764 12436
rect 4712 12393 4721 12427
rect 4721 12393 4755 12427
rect 4755 12393 4764 12427
rect 4712 12384 4764 12393
rect 4804 12384 4856 12436
rect 7104 12427 7156 12436
rect 7104 12393 7113 12427
rect 7113 12393 7147 12427
rect 7147 12393 7156 12427
rect 7104 12384 7156 12393
rect 7656 12384 7708 12436
rect 8668 12384 8720 12436
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 9680 12427 9732 12436
rect 9680 12393 9689 12427
rect 9689 12393 9723 12427
rect 9723 12393 9732 12427
rect 9680 12384 9732 12393
rect 2872 12316 2924 12368
rect 3608 12248 3660 12300
rect 2872 12223 2924 12232
rect 2872 12189 2881 12223
rect 2881 12189 2915 12223
rect 2915 12189 2924 12223
rect 2872 12180 2924 12189
rect 3424 12223 3476 12232
rect 3424 12189 3434 12223
rect 3434 12189 3476 12223
rect 3424 12180 3476 12189
rect 4528 12180 4580 12232
rect 4804 12223 4856 12232
rect 3884 12112 3936 12164
rect 3976 12112 4028 12164
rect 4804 12189 4813 12223
rect 4813 12189 4847 12223
rect 4847 12189 4856 12223
rect 4804 12180 4856 12189
rect 4988 12248 5040 12300
rect 5172 12291 5224 12300
rect 5172 12257 5181 12291
rect 5181 12257 5215 12291
rect 5215 12257 5224 12291
rect 5816 12359 5868 12368
rect 5816 12325 5825 12359
rect 5825 12325 5859 12359
rect 5859 12325 5868 12359
rect 5816 12316 5868 12325
rect 6828 12316 6880 12368
rect 10784 12316 10836 12368
rect 5172 12248 5224 12257
rect 6736 12291 6788 12300
rect 6736 12257 6745 12291
rect 6745 12257 6779 12291
rect 6779 12257 6788 12291
rect 6736 12248 6788 12257
rect 2964 12044 3016 12096
rect 5080 12112 5132 12164
rect 5540 12112 5592 12164
rect 6828 12112 6880 12164
rect 7932 12180 7984 12232
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 9312 12044 9364 12096
rect 9588 12044 9640 12096
rect 9956 12044 10008 12096
rect 11520 12044 11572 12096
rect 3036 11942 3088 11994
rect 3100 11942 3152 11994
rect 3164 11942 3216 11994
rect 3228 11942 3280 11994
rect 3292 11942 3344 11994
rect 5888 11942 5940 11994
rect 5952 11942 6004 11994
rect 6016 11942 6068 11994
rect 6080 11942 6132 11994
rect 6144 11942 6196 11994
rect 8740 11942 8792 11994
rect 8804 11942 8856 11994
rect 8868 11942 8920 11994
rect 8932 11942 8984 11994
rect 8996 11942 9048 11994
rect 11592 11942 11644 11994
rect 11656 11942 11708 11994
rect 11720 11942 11772 11994
rect 11784 11942 11836 11994
rect 11848 11942 11900 11994
rect 2780 11840 2832 11892
rect 2872 11840 2924 11892
rect 3884 11883 3936 11892
rect 3884 11849 3893 11883
rect 3893 11849 3927 11883
rect 3927 11849 3936 11883
rect 3884 11840 3936 11849
rect 4620 11840 4672 11892
rect 4896 11840 4948 11892
rect 5172 11840 5224 11892
rect 7656 11883 7708 11892
rect 7656 11849 7665 11883
rect 7665 11849 7699 11883
rect 7699 11849 7708 11883
rect 7656 11840 7708 11849
rect 8668 11840 8720 11892
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 9588 11840 9640 11892
rect 5264 11772 5316 11824
rect 1032 11704 1084 11756
rect 2964 11704 3016 11756
rect 3424 11704 3476 11756
rect 3700 11679 3752 11688
rect 3700 11645 3709 11679
rect 3709 11645 3743 11679
rect 3743 11645 3752 11679
rect 3700 11636 3752 11645
rect 3976 11747 4028 11756
rect 3976 11713 3985 11747
rect 3985 11713 4019 11747
rect 4019 11713 4028 11747
rect 3976 11704 4028 11713
rect 4068 11704 4120 11756
rect 5540 11704 5592 11756
rect 6644 11704 6696 11756
rect 7288 11747 7340 11756
rect 7288 11713 7297 11747
rect 7297 11713 7331 11747
rect 7331 11713 7340 11747
rect 7288 11704 7340 11713
rect 2872 11568 2924 11620
rect 5724 11636 5776 11688
rect 7840 11704 7892 11756
rect 7564 11636 7616 11688
rect 8484 11636 8536 11688
rect 9588 11704 9640 11756
rect 6276 11568 6328 11620
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 11520 11772 11572 11824
rect 2964 11500 3016 11552
rect 4344 11500 4396 11552
rect 4804 11500 4856 11552
rect 5632 11500 5684 11552
rect 7288 11500 7340 11552
rect 7748 11500 7800 11552
rect 8576 11500 8628 11552
rect 10600 11500 10652 11552
rect 2376 11398 2428 11450
rect 2440 11398 2492 11450
rect 2504 11398 2556 11450
rect 2568 11398 2620 11450
rect 2632 11398 2684 11450
rect 5228 11398 5280 11450
rect 5292 11398 5344 11450
rect 5356 11398 5408 11450
rect 5420 11398 5472 11450
rect 5484 11398 5536 11450
rect 8080 11398 8132 11450
rect 8144 11398 8196 11450
rect 8208 11398 8260 11450
rect 8272 11398 8324 11450
rect 8336 11398 8388 11450
rect 10932 11398 10984 11450
rect 10996 11398 11048 11450
rect 11060 11398 11112 11450
rect 11124 11398 11176 11450
rect 11188 11398 11240 11450
rect 1676 11296 1728 11348
rect 2412 11296 2464 11348
rect 2872 11296 2924 11348
rect 2964 11228 3016 11280
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2596 11067 2648 11076
rect 2596 11033 2605 11067
rect 2605 11033 2639 11067
rect 2639 11033 2648 11067
rect 2596 11024 2648 11033
rect 2780 11067 2832 11076
rect 2780 11033 2821 11067
rect 2821 11033 2832 11067
rect 3424 11296 3476 11348
rect 3700 11296 3752 11348
rect 3976 11296 4028 11348
rect 4528 11296 4580 11348
rect 5080 11296 5132 11348
rect 5724 11339 5776 11348
rect 5724 11305 5733 11339
rect 5733 11305 5767 11339
rect 5767 11305 5776 11339
rect 5724 11296 5776 11305
rect 7012 11296 7064 11348
rect 4344 11228 4396 11280
rect 3884 11160 3936 11212
rect 4068 11160 4120 11212
rect 6644 11271 6696 11280
rect 6644 11237 6653 11271
rect 6653 11237 6687 11271
rect 6687 11237 6696 11271
rect 6644 11228 6696 11237
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 10692 11296 10744 11348
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 2780 11024 2832 11033
rect 3148 11024 3200 11076
rect 4068 11067 4120 11076
rect 4068 11033 4077 11067
rect 4077 11033 4111 11067
rect 4111 11033 4120 11067
rect 4068 11024 4120 11033
rect 4160 11067 4212 11076
rect 4160 11033 4169 11067
rect 4169 11033 4203 11067
rect 4203 11033 4212 11067
rect 4160 11024 4212 11033
rect 2964 10999 3016 11008
rect 2964 10965 2973 10999
rect 2973 10965 3007 10999
rect 3007 10965 3016 10999
rect 2964 10956 3016 10965
rect 4712 11092 4764 11144
rect 4896 11067 4948 11076
rect 4896 11033 4905 11067
rect 4905 11033 4939 11067
rect 4939 11033 4948 11067
rect 4896 11024 4948 11033
rect 5080 10956 5132 11008
rect 5632 11024 5684 11076
rect 6276 11067 6328 11076
rect 6276 11033 6285 11067
rect 6285 11033 6319 11067
rect 6319 11033 6328 11067
rect 6276 11024 6328 11033
rect 7196 11160 7248 11212
rect 7564 11203 7616 11212
rect 7564 11169 7573 11203
rect 7573 11169 7607 11203
rect 7607 11169 7616 11203
rect 7564 11160 7616 11169
rect 11520 11203 11572 11212
rect 11520 11169 11529 11203
rect 11529 11169 11563 11203
rect 11563 11169 11572 11203
rect 11520 11160 11572 11169
rect 7656 11135 7708 11144
rect 7656 11101 7665 11135
rect 7665 11101 7699 11135
rect 7699 11101 7708 11135
rect 7656 11092 7708 11101
rect 6828 11024 6880 11076
rect 7840 11135 7892 11144
rect 7840 11101 7849 11135
rect 7849 11101 7883 11135
rect 7883 11101 7892 11135
rect 7840 11092 7892 11101
rect 7932 11092 7984 11144
rect 8484 11092 8536 11144
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 10784 11092 10836 11144
rect 6920 10956 6972 11008
rect 7380 10999 7432 11008
rect 7380 10965 7389 10999
rect 7389 10965 7423 10999
rect 7423 10965 7432 10999
rect 7380 10956 7432 10965
rect 10876 11024 10928 11076
rect 3036 10854 3088 10906
rect 3100 10854 3152 10906
rect 3164 10854 3216 10906
rect 3228 10854 3280 10906
rect 3292 10854 3344 10906
rect 5888 10854 5940 10906
rect 5952 10854 6004 10906
rect 6016 10854 6068 10906
rect 6080 10854 6132 10906
rect 6144 10854 6196 10906
rect 8740 10854 8792 10906
rect 8804 10854 8856 10906
rect 8868 10854 8920 10906
rect 8932 10854 8984 10906
rect 8996 10854 9048 10906
rect 11592 10854 11644 10906
rect 11656 10854 11708 10906
rect 11720 10854 11772 10906
rect 11784 10854 11836 10906
rect 11848 10854 11900 10906
rect 4344 10795 4396 10804
rect 4344 10761 4353 10795
rect 4353 10761 4387 10795
rect 4387 10761 4396 10795
rect 4344 10752 4396 10761
rect 4896 10752 4948 10804
rect 5632 10752 5684 10804
rect 7196 10752 7248 10804
rect 1676 10684 1728 10736
rect 2596 10684 2648 10736
rect 6276 10684 6328 10736
rect 10876 10684 10928 10736
rect 1952 10616 2004 10668
rect 2412 10659 2464 10668
rect 2412 10625 2421 10659
rect 2421 10625 2455 10659
rect 2455 10625 2464 10659
rect 2412 10616 2464 10625
rect 2780 10616 2832 10668
rect 2964 10616 3016 10668
rect 3608 10548 3660 10600
rect 4160 10616 4212 10668
rect 4620 10616 4672 10668
rect 7012 10616 7064 10668
rect 10232 10616 10284 10668
rect 10692 10616 10744 10668
rect 4068 10548 4120 10600
rect 4804 10480 4856 10532
rect 10784 10548 10836 10600
rect 2964 10412 3016 10464
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 5080 10455 5132 10464
rect 5080 10421 5089 10455
rect 5089 10421 5123 10455
rect 5123 10421 5132 10455
rect 5080 10412 5132 10421
rect 6920 10412 6972 10464
rect 10784 10412 10836 10464
rect 11980 10412 12032 10464
rect 2376 10310 2428 10362
rect 2440 10310 2492 10362
rect 2504 10310 2556 10362
rect 2568 10310 2620 10362
rect 2632 10310 2684 10362
rect 5228 10310 5280 10362
rect 5292 10310 5344 10362
rect 5356 10310 5408 10362
rect 5420 10310 5472 10362
rect 5484 10310 5536 10362
rect 8080 10310 8132 10362
rect 8144 10310 8196 10362
rect 8208 10310 8260 10362
rect 8272 10310 8324 10362
rect 8336 10310 8388 10362
rect 10932 10310 10984 10362
rect 10996 10310 11048 10362
rect 11060 10310 11112 10362
rect 11124 10310 11176 10362
rect 11188 10310 11240 10362
rect 4712 10208 4764 10260
rect 10232 10208 10284 10260
rect 2872 10140 2924 10192
rect 7104 10183 7156 10192
rect 7104 10149 7113 10183
rect 7113 10149 7147 10183
rect 7147 10149 7156 10183
rect 7104 10140 7156 10149
rect 6828 10047 6880 10056
rect 6828 10013 6837 10047
rect 6837 10013 6871 10047
rect 6871 10013 6880 10047
rect 6828 10004 6880 10013
rect 7380 10004 7432 10056
rect 10232 10047 10284 10056
rect 10232 10013 10241 10047
rect 10241 10013 10275 10047
rect 10275 10013 10284 10047
rect 10232 10004 10284 10013
rect 11428 10072 11480 10124
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 2964 9979 3016 9988
rect 2964 9945 2973 9979
rect 2973 9945 3007 9979
rect 3007 9945 3016 9979
rect 2964 9936 3016 9945
rect 3424 9868 3476 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7656 9868 7708 9920
rect 11336 9868 11388 9920
rect 3036 9766 3088 9818
rect 3100 9766 3152 9818
rect 3164 9766 3216 9818
rect 3228 9766 3280 9818
rect 3292 9766 3344 9818
rect 5888 9766 5940 9818
rect 5952 9766 6004 9818
rect 6016 9766 6068 9818
rect 6080 9766 6132 9818
rect 6144 9766 6196 9818
rect 8740 9766 8792 9818
rect 8804 9766 8856 9818
rect 8868 9766 8920 9818
rect 8932 9766 8984 9818
rect 8996 9766 9048 9818
rect 11592 9766 11644 9818
rect 11656 9766 11708 9818
rect 11720 9766 11772 9818
rect 11784 9766 11836 9818
rect 11848 9766 11900 9818
rect 4160 9664 4212 9716
rect 6828 9664 6880 9716
rect 2872 9596 2924 9648
rect 4804 9639 4856 9648
rect 4804 9605 4813 9639
rect 4813 9605 4847 9639
rect 4847 9605 4856 9639
rect 4804 9596 4856 9605
rect 7196 9707 7248 9716
rect 7196 9673 7205 9707
rect 7205 9673 7239 9707
rect 7239 9673 7248 9707
rect 7196 9664 7248 9673
rect 2136 9559 2148 9580
rect 2148 9559 2182 9580
rect 2182 9559 2188 9580
rect 2136 9528 2188 9559
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3424 9528 3476 9580
rect 2228 9460 2280 9512
rect 2596 9503 2648 9512
rect 2596 9469 2605 9503
rect 2605 9469 2639 9503
rect 2639 9469 2648 9503
rect 2596 9460 2648 9469
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 3976 9460 4028 9512
rect 5724 9528 5776 9580
rect 7104 9528 7156 9580
rect 7380 9639 7432 9648
rect 7380 9605 7389 9639
rect 7389 9605 7423 9639
rect 7423 9605 7432 9639
rect 7380 9596 7432 9605
rect 7748 9596 7800 9648
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 3700 9392 3752 9444
rect 4804 9392 4856 9444
rect 6920 9503 6972 9512
rect 6920 9469 6929 9503
rect 6929 9469 6963 9503
rect 6963 9469 6972 9503
rect 6920 9460 6972 9469
rect 8668 9528 8720 9580
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 5816 9367 5868 9376
rect 5816 9333 5825 9367
rect 5825 9333 5859 9367
rect 5859 9333 5868 9367
rect 5816 9324 5868 9333
rect 5908 9324 5960 9376
rect 6092 9367 6144 9376
rect 6092 9333 6101 9367
rect 6101 9333 6135 9367
rect 6135 9333 6144 9367
rect 6092 9324 6144 9333
rect 6736 9324 6788 9376
rect 6828 9324 6880 9376
rect 9128 9392 9180 9444
rect 8484 9324 8536 9376
rect 2376 9222 2428 9274
rect 2440 9222 2492 9274
rect 2504 9222 2556 9274
rect 2568 9222 2620 9274
rect 2632 9222 2684 9274
rect 5228 9222 5280 9274
rect 5292 9222 5344 9274
rect 5356 9222 5408 9274
rect 5420 9222 5472 9274
rect 5484 9222 5536 9274
rect 8080 9222 8132 9274
rect 8144 9222 8196 9274
rect 8208 9222 8260 9274
rect 8272 9222 8324 9274
rect 8336 9222 8388 9274
rect 10932 9222 10984 9274
rect 10996 9222 11048 9274
rect 11060 9222 11112 9274
rect 11124 9222 11176 9274
rect 11188 9222 11240 9274
rect 2136 9052 2188 9104
rect 2412 9052 2464 9104
rect 1492 9027 1544 9036
rect 1492 8993 1501 9027
rect 1501 8993 1535 9027
rect 1535 8993 1544 9027
rect 1492 8984 1544 8993
rect 2780 9052 2832 9104
rect 2136 8916 2188 8968
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 2964 8984 3016 9036
rect 2228 8780 2280 8832
rect 2320 8780 2372 8832
rect 3516 9052 3568 9104
rect 4252 9163 4304 9172
rect 4252 9129 4261 9163
rect 4261 9129 4295 9163
rect 4295 9129 4304 9163
rect 4252 9120 4304 9129
rect 5816 9120 5868 9172
rect 10232 9120 10284 9172
rect 4160 8984 4212 9036
rect 4988 9095 5040 9104
rect 4988 9061 4997 9095
rect 4997 9061 5031 9095
rect 5031 9061 5040 9095
rect 4988 9052 5040 9061
rect 6092 9052 6144 9104
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 3608 8959 3660 8968
rect 3608 8925 3617 8959
rect 3617 8925 3651 8959
rect 3651 8925 3660 8959
rect 3608 8916 3660 8925
rect 3792 8959 3844 8968
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 4528 8916 4580 8968
rect 5264 8916 5316 8968
rect 6276 8984 6328 9036
rect 8576 9052 8628 9104
rect 10324 9052 10376 9104
rect 7564 8984 7616 9036
rect 7748 8984 7800 9036
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 7380 8916 7432 8968
rect 8024 8916 8076 8968
rect 9404 8984 9456 9036
rect 8300 8959 8352 8968
rect 8300 8925 8309 8959
rect 8309 8925 8343 8959
rect 8343 8925 8352 8959
rect 8300 8916 8352 8925
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 9772 8959 9824 8968
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 10692 9027 10744 9036
rect 10692 8993 10701 9027
rect 10701 8993 10735 9027
rect 10735 8993 10744 9027
rect 10692 8984 10744 8993
rect 7656 8848 7708 8900
rect 8116 8891 8168 8900
rect 8116 8857 8125 8891
rect 8125 8857 8159 8891
rect 8159 8857 8168 8891
rect 8116 8848 8168 8857
rect 11336 8916 11388 8968
rect 10324 8891 10376 8900
rect 10324 8857 10333 8891
rect 10333 8857 10367 8891
rect 10367 8857 10376 8891
rect 10324 8848 10376 8857
rect 10508 8848 10560 8900
rect 11244 8848 11296 8900
rect 9588 8780 9640 8832
rect 9772 8780 9824 8832
rect 11520 8780 11572 8832
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 3036 8678 3088 8730
rect 3100 8678 3152 8730
rect 3164 8678 3216 8730
rect 3228 8678 3280 8730
rect 3292 8678 3344 8730
rect 5888 8678 5940 8730
rect 5952 8678 6004 8730
rect 6016 8678 6068 8730
rect 6080 8678 6132 8730
rect 6144 8678 6196 8730
rect 8740 8678 8792 8730
rect 8804 8678 8856 8730
rect 8868 8678 8920 8730
rect 8932 8678 8984 8730
rect 8996 8678 9048 8730
rect 11592 8678 11644 8730
rect 11656 8678 11708 8730
rect 11720 8678 11772 8730
rect 11784 8678 11836 8730
rect 11848 8678 11900 8730
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 2136 8576 2188 8585
rect 1676 8551 1728 8560
rect 1676 8517 1685 8551
rect 1685 8517 1719 8551
rect 1719 8517 1728 8551
rect 1676 8508 1728 8517
rect 2136 8440 2188 8492
rect 3332 8576 3384 8628
rect 3424 8576 3476 8628
rect 3792 8576 3844 8628
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 4160 8619 4212 8628
rect 4160 8585 4169 8619
rect 4169 8585 4203 8619
rect 4203 8585 4212 8619
rect 4160 8576 4212 8585
rect 2412 8508 2464 8560
rect 5632 8576 5684 8628
rect 3148 8483 3200 8492
rect 3148 8449 3157 8483
rect 3157 8449 3191 8483
rect 3191 8449 3200 8483
rect 3148 8440 3200 8449
rect 2228 8372 2280 8424
rect 3516 8440 3568 8492
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 4068 8440 4120 8492
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 3976 8372 4028 8424
rect 4528 8304 4580 8356
rect 5264 8551 5316 8560
rect 5264 8517 5273 8551
rect 5273 8517 5307 8551
rect 5307 8517 5316 8551
rect 5264 8508 5316 8517
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 7104 8576 7156 8628
rect 8024 8619 8076 8628
rect 8024 8585 8033 8619
rect 8033 8585 8067 8619
rect 8067 8585 8076 8619
rect 8024 8576 8076 8585
rect 9588 8576 9640 8628
rect 11336 8619 11388 8628
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 8116 8508 8168 8560
rect 6828 8372 6880 8424
rect 6368 8304 6420 8356
rect 8484 8440 8536 8492
rect 7748 8304 7800 8356
rect 9128 8440 9180 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 10324 8440 10376 8492
rect 9864 8372 9916 8424
rect 10692 8440 10744 8492
rect 10784 8372 10836 8424
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 1860 8279 1912 8288
rect 1860 8245 1869 8279
rect 1869 8245 1903 8279
rect 1903 8245 1912 8279
rect 1860 8236 1912 8245
rect 2872 8236 2924 8288
rect 3608 8236 3660 8288
rect 3700 8236 3752 8288
rect 5356 8236 5408 8288
rect 5724 8236 5776 8288
rect 7196 8236 7248 8288
rect 8300 8236 8352 8288
rect 10324 8304 10376 8356
rect 11336 8304 11388 8356
rect 10508 8236 10560 8288
rect 2376 8134 2428 8186
rect 2440 8134 2492 8186
rect 2504 8134 2556 8186
rect 2568 8134 2620 8186
rect 2632 8134 2684 8186
rect 5228 8134 5280 8186
rect 5292 8134 5344 8186
rect 5356 8134 5408 8186
rect 5420 8134 5472 8186
rect 5484 8134 5536 8186
rect 8080 8134 8132 8186
rect 8144 8134 8196 8186
rect 8208 8134 8260 8186
rect 8272 8134 8324 8186
rect 8336 8134 8388 8186
rect 10932 8134 10984 8186
rect 10996 8134 11048 8186
rect 11060 8134 11112 8186
rect 11124 8134 11176 8186
rect 11188 8134 11240 8186
rect 1308 8032 1360 8084
rect 2044 8032 2096 8084
rect 2228 8032 2280 8084
rect 3516 8032 3568 8084
rect 4436 8032 4488 8084
rect 5908 8032 5960 8084
rect 9496 8032 9548 8084
rect 10784 8032 10836 8084
rect 1492 8007 1544 8016
rect 1492 7973 1501 8007
rect 1501 7973 1535 8007
rect 1535 7973 1544 8007
rect 1492 7964 1544 7973
rect 1676 7964 1728 8016
rect 2504 7964 2556 8016
rect 2872 7964 2924 8016
rect 10968 8007 11020 8016
rect 10968 7973 10977 8007
rect 10977 7973 11011 8007
rect 11011 7973 11020 8007
rect 10968 7964 11020 7973
rect 4988 7896 5040 7948
rect 6552 7896 6604 7948
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2136 7828 2188 7880
rect 2504 7828 2556 7880
rect 2688 7871 2740 7880
rect 2688 7837 2697 7871
rect 2697 7837 2731 7871
rect 2731 7837 2740 7871
rect 2688 7828 2740 7837
rect 1860 7760 1912 7812
rect 3884 7828 3936 7880
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 5080 7828 5132 7880
rect 5632 7828 5684 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 7104 7828 7156 7880
rect 8116 7828 8168 7880
rect 3976 7760 4028 7812
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 11796 7871 11848 7880
rect 11796 7837 11805 7871
rect 11805 7837 11839 7871
rect 11839 7837 11848 7871
rect 11796 7828 11848 7837
rect 10508 7760 10560 7812
rect 2872 7692 2924 7744
rect 5080 7692 5132 7744
rect 7932 7692 7984 7744
rect 11428 7735 11480 7744
rect 11428 7701 11437 7735
rect 11437 7701 11471 7735
rect 11471 7701 11480 7735
rect 11428 7692 11480 7701
rect 3036 7590 3088 7642
rect 3100 7590 3152 7642
rect 3164 7590 3216 7642
rect 3228 7590 3280 7642
rect 3292 7590 3344 7642
rect 5888 7590 5940 7642
rect 5952 7590 6004 7642
rect 6016 7590 6068 7642
rect 6080 7590 6132 7642
rect 6144 7590 6196 7642
rect 8740 7590 8792 7642
rect 8804 7590 8856 7642
rect 8868 7590 8920 7642
rect 8932 7590 8984 7642
rect 8996 7590 9048 7642
rect 11592 7590 11644 7642
rect 11656 7590 11708 7642
rect 11720 7590 11772 7642
rect 11784 7590 11836 7642
rect 11848 7590 11900 7642
rect 940 7420 992 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2872 7463 2924 7472
rect 2872 7429 2881 7463
rect 2881 7429 2915 7463
rect 2915 7429 2924 7463
rect 2872 7420 2924 7429
rect 3976 7420 4028 7472
rect 6552 7531 6604 7540
rect 6552 7497 6561 7531
rect 6561 7497 6595 7531
rect 6595 7497 6604 7531
rect 6552 7488 6604 7497
rect 10416 7488 10468 7540
rect 1952 7352 2004 7404
rect 2688 7284 2740 7336
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 3792 7352 3844 7404
rect 10508 7463 10560 7472
rect 10508 7429 10517 7463
rect 10517 7429 10551 7463
rect 10551 7429 10560 7463
rect 10508 7420 10560 7429
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 6736 7352 6788 7404
rect 2136 7216 2188 7268
rect 3884 7216 3936 7268
rect 7012 7284 7064 7336
rect 7932 7395 7984 7404
rect 7932 7361 7941 7395
rect 7941 7361 7975 7395
rect 7975 7361 7984 7395
rect 7932 7352 7984 7361
rect 8024 7352 8076 7404
rect 10140 7352 10192 7404
rect 11520 7488 11572 7540
rect 10692 7395 10744 7404
rect 10692 7361 10701 7395
rect 10701 7361 10735 7395
rect 10735 7361 10744 7395
rect 10968 7395 11020 7404
rect 10692 7352 10744 7361
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 11428 7352 11480 7404
rect 11520 7395 11572 7404
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 11980 7352 12032 7404
rect 7840 7284 7892 7336
rect 8116 7327 8168 7336
rect 8116 7293 8125 7327
rect 8125 7293 8159 7327
rect 8159 7293 8168 7327
rect 8116 7284 8168 7293
rect 11336 7284 11388 7336
rect 7472 7216 7524 7268
rect 10876 7216 10928 7268
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 2228 7148 2280 7200
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 8484 7148 8536 7200
rect 9956 7148 10008 7200
rect 2376 7046 2428 7098
rect 2440 7046 2492 7098
rect 2504 7046 2556 7098
rect 2568 7046 2620 7098
rect 2632 7046 2684 7098
rect 5228 7046 5280 7098
rect 5292 7046 5344 7098
rect 5356 7046 5408 7098
rect 5420 7046 5472 7098
rect 5484 7046 5536 7098
rect 8080 7046 8132 7098
rect 8144 7046 8196 7098
rect 8208 7046 8260 7098
rect 8272 7046 8324 7098
rect 8336 7046 8388 7098
rect 10932 7046 10984 7098
rect 10996 7046 11048 7098
rect 11060 7046 11112 7098
rect 11124 7046 11176 7098
rect 11188 7046 11240 7098
rect 1676 6944 1728 6996
rect 7472 6987 7524 6996
rect 7472 6953 7481 6987
rect 7481 6953 7515 6987
rect 7515 6953 7524 6987
rect 7472 6944 7524 6953
rect 5356 6876 5408 6928
rect 7012 6876 7064 6928
rect 10048 6876 10100 6928
rect 11980 6876 12032 6928
rect 2872 6808 2924 6860
rect 2596 6740 2648 6792
rect 2136 6672 2188 6724
rect 2228 6604 2280 6656
rect 2964 6604 3016 6656
rect 3332 6740 3384 6792
rect 4896 6740 4948 6792
rect 7932 6808 7984 6860
rect 3700 6672 3752 6724
rect 7196 6672 7248 6724
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 8484 6740 8536 6792
rect 10508 6808 10560 6860
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 11428 6808 11480 6860
rect 12164 6851 12216 6860
rect 12164 6817 12173 6851
rect 12173 6817 12207 6851
rect 12207 6817 12216 6851
rect 12164 6808 12216 6817
rect 11336 6740 11388 6792
rect 3792 6604 3844 6656
rect 5172 6604 5224 6656
rect 5356 6647 5408 6656
rect 5356 6613 5365 6647
rect 5365 6613 5399 6647
rect 5399 6613 5408 6647
rect 5356 6604 5408 6613
rect 6276 6604 6328 6656
rect 7472 6604 7524 6656
rect 9220 6672 9272 6724
rect 8484 6604 8536 6656
rect 9496 6604 9548 6656
rect 10968 6604 11020 6656
rect 3036 6502 3088 6554
rect 3100 6502 3152 6554
rect 3164 6502 3216 6554
rect 3228 6502 3280 6554
rect 3292 6502 3344 6554
rect 5888 6502 5940 6554
rect 5952 6502 6004 6554
rect 6016 6502 6068 6554
rect 6080 6502 6132 6554
rect 6144 6502 6196 6554
rect 8740 6502 8792 6554
rect 8804 6502 8856 6554
rect 8868 6502 8920 6554
rect 8932 6502 8984 6554
rect 8996 6502 9048 6554
rect 11592 6502 11644 6554
rect 11656 6502 11708 6554
rect 11720 6502 11772 6554
rect 11784 6502 11836 6554
rect 11848 6502 11900 6554
rect 2596 6443 2648 6452
rect 2596 6409 2605 6443
rect 2605 6409 2639 6443
rect 2639 6409 2648 6443
rect 2596 6400 2648 6409
rect 4896 6400 4948 6452
rect 2964 6332 3016 6384
rect 7104 6400 7156 6452
rect 7380 6400 7432 6452
rect 848 6264 900 6316
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 2780 6264 2832 6273
rect 2872 6239 2924 6248
rect 2872 6205 2881 6239
rect 2881 6205 2915 6239
rect 2915 6205 2924 6239
rect 2872 6196 2924 6205
rect 3148 6196 3200 6248
rect 4068 6307 4120 6316
rect 4068 6273 4077 6307
rect 4077 6273 4111 6307
rect 4111 6273 4120 6307
rect 4068 6264 4120 6273
rect 4712 6264 4764 6316
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 6368 6332 6420 6384
rect 2780 6060 2832 6112
rect 3792 6171 3844 6180
rect 3792 6137 3801 6171
rect 3801 6137 3835 6171
rect 3835 6137 3844 6171
rect 3792 6128 3844 6137
rect 4988 6239 5040 6248
rect 4988 6205 4997 6239
rect 4997 6205 5031 6239
rect 5031 6205 5040 6239
rect 4988 6196 5040 6205
rect 5816 6307 5868 6316
rect 5816 6273 5825 6307
rect 5825 6273 5859 6307
rect 5859 6273 5868 6307
rect 5816 6264 5868 6273
rect 7104 6264 7156 6316
rect 5448 6128 5500 6180
rect 7380 6196 7432 6248
rect 4804 6060 4856 6112
rect 5632 6060 5684 6112
rect 8484 6307 8536 6316
rect 8484 6273 8493 6307
rect 8493 6273 8527 6307
rect 8527 6273 8536 6307
rect 8484 6264 8536 6273
rect 9496 6332 9548 6384
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 8576 6196 8628 6248
rect 10232 6264 10284 6316
rect 10784 6375 10836 6384
rect 10784 6341 10793 6375
rect 10793 6341 10827 6375
rect 10827 6341 10836 6375
rect 10784 6332 10836 6341
rect 10968 6443 11020 6452
rect 10968 6409 10977 6443
rect 10977 6409 11011 6443
rect 11011 6409 11020 6443
rect 10968 6400 11020 6409
rect 11520 6400 11572 6452
rect 11980 6375 12032 6384
rect 11980 6341 11989 6375
rect 11989 6341 12023 6375
rect 12023 6341 12032 6375
rect 11980 6332 12032 6341
rect 10416 6239 10468 6248
rect 10416 6205 10425 6239
rect 10425 6205 10459 6239
rect 10459 6205 10468 6239
rect 10416 6196 10468 6205
rect 9220 6171 9272 6180
rect 9220 6137 9229 6171
rect 9229 6137 9263 6171
rect 9263 6137 9272 6171
rect 9220 6128 9272 6137
rect 11336 6128 11388 6180
rect 11612 6171 11664 6180
rect 11612 6137 11621 6171
rect 11621 6137 11655 6171
rect 11655 6137 11664 6171
rect 11612 6128 11664 6137
rect 9772 6103 9824 6112
rect 9772 6069 9781 6103
rect 9781 6069 9815 6103
rect 9815 6069 9824 6103
rect 9772 6060 9824 6069
rect 11428 6060 11480 6112
rect 2376 5958 2428 6010
rect 2440 5958 2492 6010
rect 2504 5958 2556 6010
rect 2568 5958 2620 6010
rect 2632 5958 2684 6010
rect 5228 5958 5280 6010
rect 5292 5958 5344 6010
rect 5356 5958 5408 6010
rect 5420 5958 5472 6010
rect 5484 5958 5536 6010
rect 8080 5958 8132 6010
rect 8144 5958 8196 6010
rect 8208 5958 8260 6010
rect 8272 5958 8324 6010
rect 8336 5958 8388 6010
rect 10932 5958 10984 6010
rect 10996 5958 11048 6010
rect 11060 5958 11112 6010
rect 11124 5958 11176 6010
rect 11188 5958 11240 6010
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 3424 5856 3476 5908
rect 4712 5856 4764 5908
rect 3700 5788 3752 5840
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 5724 5856 5776 5908
rect 6000 5856 6052 5908
rect 6368 5856 6420 5908
rect 9036 5856 9088 5908
rect 10508 5856 10560 5908
rect 3516 5720 3568 5772
rect 1492 5627 1544 5636
rect 1492 5593 1501 5627
rect 1501 5593 1535 5627
rect 1535 5593 1544 5627
rect 1492 5584 1544 5593
rect 2228 5627 2280 5636
rect 2228 5593 2237 5627
rect 2237 5593 2271 5627
rect 2271 5593 2280 5627
rect 2228 5584 2280 5593
rect 2688 5652 2740 5704
rect 2872 5652 2924 5704
rect 10416 5788 10468 5840
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 4068 5652 4120 5704
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 4896 5652 4948 5704
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 4528 5584 4580 5636
rect 2872 5516 2924 5568
rect 3424 5516 3476 5568
rect 4344 5516 4396 5568
rect 5816 5652 5868 5704
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 7104 5652 7156 5704
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 7380 5652 7432 5704
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 9220 5720 9272 5772
rect 9772 5720 9824 5772
rect 8576 5652 8628 5704
rect 10232 5652 10284 5704
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 5172 5516 5224 5568
rect 5632 5516 5684 5568
rect 6276 5516 6328 5568
rect 7748 5559 7800 5568
rect 7748 5525 7757 5559
rect 7757 5525 7791 5559
rect 7791 5525 7800 5559
rect 7748 5516 7800 5525
rect 8668 5584 8720 5636
rect 10140 5584 10192 5636
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 11336 5720 11388 5772
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 10692 5516 10744 5568
rect 3036 5414 3088 5466
rect 3100 5414 3152 5466
rect 3164 5414 3216 5466
rect 3228 5414 3280 5466
rect 3292 5414 3344 5466
rect 5888 5414 5940 5466
rect 5952 5414 6004 5466
rect 6016 5414 6068 5466
rect 6080 5414 6132 5466
rect 6144 5414 6196 5466
rect 8740 5414 8792 5466
rect 8804 5414 8856 5466
rect 8868 5414 8920 5466
rect 8932 5414 8984 5466
rect 8996 5414 9048 5466
rect 11592 5414 11644 5466
rect 11656 5414 11708 5466
rect 11720 5414 11772 5466
rect 11784 5414 11836 5466
rect 11848 5414 11900 5466
rect 4068 5312 4120 5364
rect 7288 5312 7340 5364
rect 10508 5312 10560 5364
rect 12072 5355 12124 5364
rect 12072 5321 12081 5355
rect 12081 5321 12115 5355
rect 12115 5321 12124 5355
rect 12072 5312 12124 5321
rect 2228 5244 2280 5296
rect 848 5176 900 5228
rect 2780 5176 2832 5228
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 4436 5244 4488 5296
rect 5080 5244 5132 5296
rect 8576 5244 8628 5296
rect 11428 5244 11480 5296
rect 4804 5176 4856 5228
rect 7104 5176 7156 5228
rect 7932 5176 7984 5228
rect 9956 5176 10008 5228
rect 10140 5176 10192 5228
rect 2044 5108 2096 5160
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 7196 5108 7248 5160
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 7840 5108 7892 5160
rect 8484 5151 8536 5160
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 2376 4870 2428 4922
rect 2440 4870 2492 4922
rect 2504 4870 2556 4922
rect 2568 4870 2620 4922
rect 2632 4870 2684 4922
rect 5228 4870 5280 4922
rect 5292 4870 5344 4922
rect 5356 4870 5408 4922
rect 5420 4870 5472 4922
rect 5484 4870 5536 4922
rect 8080 4870 8132 4922
rect 8144 4870 8196 4922
rect 8208 4870 8260 4922
rect 8272 4870 8324 4922
rect 8336 4870 8388 4922
rect 10932 4870 10984 4922
rect 10996 4870 11048 4922
rect 11060 4870 11112 4922
rect 11124 4870 11176 4922
rect 11188 4870 11240 4922
rect 2872 4768 2924 4820
rect 3240 4768 3292 4820
rect 4068 4768 4120 4820
rect 4804 4811 4856 4820
rect 4804 4777 4813 4811
rect 4813 4777 4847 4811
rect 4847 4777 4856 4811
rect 4804 4768 4856 4777
rect 7656 4768 7708 4820
rect 7840 4768 7892 4820
rect 8484 4768 8536 4820
rect 4436 4632 4488 4684
rect 2228 4564 2280 4616
rect 3516 4564 3568 4616
rect 4160 4564 4212 4616
rect 4988 4607 5040 4616
rect 4988 4573 4997 4607
rect 4997 4573 5031 4607
rect 5031 4573 5040 4607
rect 4988 4564 5040 4573
rect 5080 4564 5132 4616
rect 6368 4564 6420 4616
rect 5632 4428 5684 4480
rect 7104 4496 7156 4548
rect 7932 4607 7984 4616
rect 7932 4573 7941 4607
rect 7941 4573 7975 4607
rect 7975 4573 7984 4607
rect 7932 4564 7984 4573
rect 8300 4564 8352 4616
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 10692 4811 10744 4820
rect 10692 4777 10701 4811
rect 10701 4777 10735 4811
rect 10735 4777 10744 4811
rect 10692 4768 10744 4777
rect 10324 4700 10376 4752
rect 11980 4768 12032 4820
rect 10416 4632 10468 4684
rect 8576 4496 8628 4548
rect 9404 4564 9456 4616
rect 9956 4564 10008 4616
rect 10968 4632 11020 4684
rect 11520 4496 11572 4548
rect 10232 4428 10284 4480
rect 11152 4471 11204 4480
rect 11152 4437 11161 4471
rect 11161 4437 11195 4471
rect 11195 4437 11204 4471
rect 11152 4428 11204 4437
rect 3036 4326 3088 4378
rect 3100 4326 3152 4378
rect 3164 4326 3216 4378
rect 3228 4326 3280 4378
rect 3292 4326 3344 4378
rect 5888 4326 5940 4378
rect 5952 4326 6004 4378
rect 6016 4326 6068 4378
rect 6080 4326 6132 4378
rect 6144 4326 6196 4378
rect 8740 4326 8792 4378
rect 8804 4326 8856 4378
rect 8868 4326 8920 4378
rect 8932 4326 8984 4378
rect 8996 4326 9048 4378
rect 11592 4326 11644 4378
rect 11656 4326 11708 4378
rect 11720 4326 11772 4378
rect 11784 4326 11836 4378
rect 11848 4326 11900 4378
rect 4436 4224 4488 4276
rect 4068 4156 4120 4208
rect 4988 4156 5040 4208
rect 4344 4088 4396 4140
rect 4436 4020 4488 4072
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 4160 3927 4212 3936
rect 4160 3893 4169 3927
rect 4169 3893 4203 3927
rect 4203 3893 4212 3927
rect 4160 3884 4212 3893
rect 4344 3927 4396 3936
rect 4344 3893 4353 3927
rect 4353 3893 4387 3927
rect 4387 3893 4396 3927
rect 4344 3884 4396 3893
rect 4620 3884 4672 3936
rect 5080 4020 5132 4072
rect 5540 4224 5592 4276
rect 10232 4224 10284 4276
rect 5724 4156 5776 4208
rect 10140 4156 10192 4208
rect 6828 4088 6880 4140
rect 7748 4088 7800 4140
rect 7932 4088 7984 4140
rect 10416 4156 10468 4208
rect 10692 4156 10744 4208
rect 10324 4131 10376 4140
rect 10324 4097 10333 4131
rect 10333 4097 10367 4131
rect 10367 4097 10376 4131
rect 10324 4088 10376 4097
rect 6368 4020 6420 4072
rect 7564 4063 7616 4072
rect 7564 4029 7573 4063
rect 7573 4029 7607 4063
rect 7607 4029 7616 4063
rect 7564 4020 7616 4029
rect 10600 4088 10652 4140
rect 11152 4156 11204 4208
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 5816 3995 5868 4004
rect 5816 3961 5825 3995
rect 5825 3961 5859 3995
rect 5859 3961 5868 3995
rect 5816 3952 5868 3961
rect 10048 3952 10100 4004
rect 10416 3995 10468 4004
rect 10416 3961 10425 3995
rect 10425 3961 10459 3995
rect 10459 3961 10468 3995
rect 10416 3952 10468 3961
rect 10784 3952 10836 4004
rect 6000 3927 6052 3936
rect 6000 3893 6009 3927
rect 6009 3893 6043 3927
rect 6043 3893 6052 3927
rect 6000 3884 6052 3893
rect 8484 3884 8536 3936
rect 9220 3884 9272 3936
rect 10324 3884 10376 3936
rect 2376 3782 2428 3834
rect 2440 3782 2492 3834
rect 2504 3782 2556 3834
rect 2568 3782 2620 3834
rect 2632 3782 2684 3834
rect 5228 3782 5280 3834
rect 5292 3782 5344 3834
rect 5356 3782 5408 3834
rect 5420 3782 5472 3834
rect 5484 3782 5536 3834
rect 8080 3782 8132 3834
rect 8144 3782 8196 3834
rect 8208 3782 8260 3834
rect 8272 3782 8324 3834
rect 8336 3782 8388 3834
rect 10932 3782 10984 3834
rect 10996 3782 11048 3834
rect 11060 3782 11112 3834
rect 11124 3782 11176 3834
rect 11188 3782 11240 3834
rect 4436 3723 4488 3732
rect 4436 3689 4445 3723
rect 4445 3689 4479 3723
rect 4479 3689 4488 3723
rect 4436 3680 4488 3689
rect 4804 3680 4856 3732
rect 6000 3723 6052 3732
rect 6000 3689 6009 3723
rect 6009 3689 6043 3723
rect 6043 3689 6052 3723
rect 6000 3680 6052 3689
rect 10416 3680 10468 3732
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4344 3519 4396 3528
rect 4344 3485 4353 3519
rect 4353 3485 4387 3519
rect 4387 3485 4396 3519
rect 4344 3476 4396 3485
rect 4436 3476 4488 3528
rect 5356 3476 5408 3528
rect 5632 3612 5684 3664
rect 5724 3544 5776 3596
rect 6460 3612 6512 3664
rect 9312 3612 9364 3664
rect 9956 3612 10008 3664
rect 6920 3544 6972 3596
rect 9772 3544 9824 3596
rect 5724 3408 5776 3460
rect 5816 3408 5868 3460
rect 6276 3451 6328 3460
rect 6276 3417 6285 3451
rect 6285 3417 6319 3451
rect 6319 3417 6328 3451
rect 6276 3408 6328 3417
rect 7104 3476 7156 3528
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 7012 3408 7064 3460
rect 6552 3340 6604 3392
rect 9404 3476 9456 3528
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10324 3476 10376 3528
rect 9312 3408 9364 3460
rect 10692 3408 10744 3460
rect 3036 3238 3088 3290
rect 3100 3238 3152 3290
rect 3164 3238 3216 3290
rect 3228 3238 3280 3290
rect 3292 3238 3344 3290
rect 5888 3238 5940 3290
rect 5952 3238 6004 3290
rect 6016 3238 6068 3290
rect 6080 3238 6132 3290
rect 6144 3238 6196 3290
rect 8740 3238 8792 3290
rect 8804 3238 8856 3290
rect 8868 3238 8920 3290
rect 8932 3238 8984 3290
rect 8996 3238 9048 3290
rect 11592 3238 11644 3290
rect 11656 3238 11708 3290
rect 11720 3238 11772 3290
rect 11784 3238 11836 3290
rect 11848 3238 11900 3290
rect 5080 3136 5132 3188
rect 5724 3136 5776 3188
rect 5816 3136 5868 3188
rect 7564 3136 7616 3188
rect 9312 3136 9364 3188
rect 10048 3136 10100 3188
rect 4160 3000 4212 3052
rect 4712 3000 4764 3052
rect 5632 3000 5684 3052
rect 4344 2932 4396 2984
rect 6276 3000 6328 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 6460 2932 6512 2984
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 7932 3043 7984 3052
rect 7932 3009 7941 3043
rect 7941 3009 7975 3043
rect 7975 3009 7984 3043
rect 7932 3000 7984 3009
rect 6552 2864 6604 2916
rect 6828 2864 6880 2916
rect 9864 3068 9916 3120
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10140 2932 10192 2984
rect 10416 3000 10468 3052
rect 10600 2932 10652 2984
rect 6276 2796 6328 2848
rect 9220 2839 9272 2848
rect 9220 2805 9229 2839
rect 9229 2805 9263 2839
rect 9263 2805 9272 2839
rect 9220 2796 9272 2805
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 10048 2796 10100 2805
rect 2376 2694 2428 2746
rect 2440 2694 2492 2746
rect 2504 2694 2556 2746
rect 2568 2694 2620 2746
rect 2632 2694 2684 2746
rect 5228 2694 5280 2746
rect 5292 2694 5344 2746
rect 5356 2694 5408 2746
rect 5420 2694 5472 2746
rect 5484 2694 5536 2746
rect 8080 2694 8132 2746
rect 8144 2694 8196 2746
rect 8208 2694 8260 2746
rect 8272 2694 8324 2746
rect 8336 2694 8388 2746
rect 10932 2694 10984 2746
rect 10996 2694 11048 2746
rect 11060 2694 11112 2746
rect 11124 2694 11176 2746
rect 11188 2694 11240 2746
rect 4988 2592 5040 2644
rect 7932 2592 7984 2644
rect 10048 2592 10100 2644
rect 5172 2524 5224 2576
rect 5724 2456 5776 2508
rect 7012 2456 7064 2508
rect 9404 2499 9456 2508
rect 9404 2465 9413 2499
rect 9413 2465 9447 2499
rect 9447 2465 9456 2499
rect 9404 2456 9456 2465
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5816 2388 5868 2440
rect 7104 2388 7156 2440
rect 8484 2388 8536 2440
rect 6460 2320 6512 2372
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9680 2388 9732 2440
rect 4528 2252 4580 2304
rect 7748 2252 7800 2304
rect 8392 2252 8444 2304
rect 3036 2150 3088 2202
rect 3100 2150 3152 2202
rect 3164 2150 3216 2202
rect 3228 2150 3280 2202
rect 3292 2150 3344 2202
rect 5888 2150 5940 2202
rect 5952 2150 6004 2202
rect 6016 2150 6068 2202
rect 6080 2150 6132 2202
rect 6144 2150 6196 2202
rect 8740 2150 8792 2202
rect 8804 2150 8856 2202
rect 8868 2150 8920 2202
rect 8932 2150 8984 2202
rect 8996 2150 9048 2202
rect 11592 2150 11644 2202
rect 11656 2150 11708 2202
rect 11720 2150 11772 2202
rect 11784 2150 11836 2202
rect 11848 2150 11900 2202
<< metal2 >>
rect 4526 14990 4582 15790
rect 6458 14990 6514 15790
rect 7102 14990 7158 15790
rect 7746 14990 7802 15790
rect 2376 13628 2684 13637
rect 2376 13626 2382 13628
rect 2438 13626 2462 13628
rect 2518 13626 2542 13628
rect 2598 13626 2622 13628
rect 2678 13626 2684 13628
rect 2438 13574 2440 13626
rect 2620 13574 2622 13626
rect 2376 13572 2382 13574
rect 2438 13572 2462 13574
rect 2518 13572 2542 13574
rect 2598 13572 2622 13574
rect 2678 13572 2684 13574
rect 2376 13563 2684 13572
rect 4540 13326 4568 14990
rect 5228 13628 5536 13637
rect 5228 13626 5234 13628
rect 5290 13626 5314 13628
rect 5370 13626 5394 13628
rect 5450 13626 5474 13628
rect 5530 13626 5536 13628
rect 5290 13574 5292 13626
rect 5472 13574 5474 13626
rect 5228 13572 5234 13574
rect 5290 13572 5314 13574
rect 5370 13572 5394 13574
rect 5450 13572 5474 13574
rect 5530 13572 5536 13574
rect 5228 13563 5536 13572
rect 6472 13326 6500 14990
rect 7116 13326 7144 14990
rect 7760 13394 7788 14990
rect 8080 13628 8388 13637
rect 8080 13626 8086 13628
rect 8142 13626 8166 13628
rect 8222 13626 8246 13628
rect 8302 13626 8326 13628
rect 8382 13626 8388 13628
rect 8142 13574 8144 13626
rect 8324 13574 8326 13626
rect 8080 13572 8086 13574
rect 8142 13572 8166 13574
rect 8222 13572 8246 13574
rect 8302 13572 8326 13574
rect 8382 13572 8388 13574
rect 8080 13563 8388 13572
rect 10932 13628 11240 13637
rect 10932 13626 10938 13628
rect 10994 13626 11018 13628
rect 11074 13626 11098 13628
rect 11154 13626 11178 13628
rect 11234 13626 11240 13628
rect 10994 13574 10996 13626
rect 11176 13574 11178 13626
rect 10932 13572 10938 13574
rect 10994 13572 11018 13574
rect 11074 13572 11098 13574
rect 11154 13572 11178 13574
rect 11234 13572 11240 13574
rect 10932 13563 11240 13572
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 3036 13084 3344 13093
rect 3036 13082 3042 13084
rect 3098 13082 3122 13084
rect 3178 13082 3202 13084
rect 3258 13082 3282 13084
rect 3338 13082 3344 13084
rect 3098 13030 3100 13082
rect 3280 13030 3282 13082
rect 3036 13028 3042 13030
rect 3098 13028 3122 13030
rect 3178 13028 3202 13030
rect 3258 13028 3282 13030
rect 3338 13028 3344 13030
rect 3036 13019 3344 13028
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1032 11756 1084 11762
rect 1032 11698 1084 11704
rect 1044 11665 1072 11698
rect 1030 11656 1086 11665
rect 1030 11591 1086 11600
rect 1688 11354 1716 12582
rect 2376 12540 2684 12549
rect 2376 12538 2382 12540
rect 2438 12538 2462 12540
rect 2518 12538 2542 12540
rect 2598 12538 2622 12540
rect 2678 12538 2684 12540
rect 2438 12486 2440 12538
rect 2620 12486 2622 12538
rect 2376 12484 2382 12486
rect 2438 12484 2462 12486
rect 2518 12484 2542 12486
rect 2598 12484 2622 12486
rect 2678 12484 2684 12486
rect 2376 12475 2684 12484
rect 2872 12368 2924 12374
rect 2792 12316 2872 12322
rect 2792 12310 2924 12316
rect 2792 12294 2912 12310
rect 3608 12300 3660 12306
rect 2792 11898 2820 12294
rect 3608 12242 3660 12248
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 2884 11898 2912 12174
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2976 11762 3004 12038
rect 3036 11996 3344 12005
rect 3036 11994 3042 11996
rect 3098 11994 3122 11996
rect 3178 11994 3202 11996
rect 3258 11994 3282 11996
rect 3338 11994 3344 11996
rect 3098 11942 3100 11994
rect 3280 11942 3282 11994
rect 3036 11940 3042 11942
rect 3098 11940 3122 11942
rect 3178 11940 3202 11942
rect 3258 11940 3282 11942
rect 3338 11940 3344 11942
rect 3036 11931 3344 11940
rect 3436 11762 3464 12174
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 3424 11756 3476 11762
rect 3424 11698 3476 11704
rect 2872 11620 2924 11626
rect 2872 11562 2924 11568
rect 2376 11452 2684 11461
rect 2376 11450 2382 11452
rect 2438 11450 2462 11452
rect 2518 11450 2542 11452
rect 2598 11450 2622 11452
rect 2678 11450 2684 11452
rect 2438 11398 2440 11450
rect 2620 11398 2622 11450
rect 2376 11396 2382 11398
rect 2438 11396 2462 11398
rect 2518 11396 2542 11398
rect 2598 11396 2622 11398
rect 2678 11396 2684 11398
rect 2376 11387 2684 11396
rect 2884 11354 2912 11562
rect 2976 11558 3004 11698
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 3436 11354 3464 11698
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1676 10736 1728 10742
rect 1676 10678 1728 10684
rect 1688 9625 1716 10678
rect 2424 10674 2452 11290
rect 2964 11280 3016 11286
rect 3016 11228 3096 11234
rect 2964 11222 3096 11228
rect 2976 11206 3096 11222
rect 2596 11076 2648 11082
rect 2596 11018 2648 11024
rect 2780 11076 2832 11082
rect 3068 11064 3096 11206
rect 3148 11076 3200 11082
rect 3068 11036 3148 11064
rect 2780 11018 2832 11024
rect 3148 11018 3200 11024
rect 2608 10742 2636 11018
rect 2596 10736 2648 10742
rect 2596 10678 2648 10684
rect 2792 10674 2820 11018
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2976 10674 3004 10950
rect 3036 10908 3344 10917
rect 3036 10906 3042 10908
rect 3098 10906 3122 10908
rect 3178 10906 3202 10908
rect 3258 10906 3282 10908
rect 3338 10906 3344 10908
rect 3098 10854 3100 10906
rect 3280 10854 3282 10906
rect 3036 10852 3042 10854
rect 3098 10852 3122 10854
rect 3178 10852 3202 10854
rect 3258 10852 3282 10854
rect 3338 10852 3344 10854
rect 3036 10843 3344 10852
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 2412 10668 2464 10674
rect 2412 10610 2464 10616
rect 2780 10668 2832 10674
rect 2964 10668 3016 10674
rect 2780 10610 2832 10616
rect 2884 10628 2964 10656
rect 1674 9616 1730 9625
rect 1674 9551 1730 9560
rect 1490 9072 1546 9081
rect 1490 9007 1492 9016
rect 1544 9007 1546 9016
rect 1492 8978 1544 8984
rect 1490 8936 1546 8945
rect 1490 8871 1546 8880
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1320 8090 1348 8191
rect 1308 8084 1360 8090
rect 1308 8026 1360 8032
rect 1504 8022 1532 8871
rect 1688 8566 1716 9551
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1688 8022 1716 8502
rect 1860 8288 1912 8294
rect 1860 8230 1912 8236
rect 1492 8016 1544 8022
rect 1492 7958 1544 7964
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1872 7818 1900 8230
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 938 7576 994 7585
rect 938 7511 994 7520
rect 952 7478 980 7511
rect 940 7472 992 7478
rect 940 7414 992 7420
rect 1964 7410 1992 10610
rect 2376 10364 2684 10373
rect 2376 10362 2382 10364
rect 2438 10362 2462 10364
rect 2518 10362 2542 10364
rect 2598 10362 2622 10364
rect 2678 10362 2684 10364
rect 2438 10310 2440 10362
rect 2620 10310 2622 10362
rect 2376 10308 2382 10310
rect 2438 10308 2462 10310
rect 2518 10308 2542 10310
rect 2598 10308 2622 10310
rect 2678 10308 2684 10310
rect 2376 10299 2684 10308
rect 2884 10198 2912 10628
rect 2964 10610 3016 10616
rect 3620 10606 3648 12242
rect 4528 12232 4580 12238
rect 4526 12200 4528 12209
rect 4580 12200 4582 12209
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3976 12164 4028 12170
rect 4526 12135 4582 12144
rect 3976 12106 4028 12112
rect 3896 11898 3924 12106
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3988 11762 4016 12106
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3712 11354 3740 11630
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2872 10192 2924 10198
rect 2872 10134 2924 10140
rect 2976 9994 3004 10406
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3036 9820 3344 9829
rect 3036 9818 3042 9820
rect 3098 9818 3122 9820
rect 3178 9818 3202 9820
rect 3258 9818 3282 9820
rect 3338 9818 3344 9820
rect 3098 9766 3100 9818
rect 3280 9766 3282 9818
rect 3036 9764 3042 9766
rect 3098 9764 3122 9766
rect 3178 9764 3202 9766
rect 3258 9764 3282 9766
rect 3338 9764 3344 9766
rect 3036 9755 3344 9764
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 3146 9616 3202 9625
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 2148 9110 2176 9522
rect 2228 9512 2280 9518
rect 2596 9512 2648 9518
rect 2228 9454 2280 9460
rect 2594 9480 2596 9489
rect 2648 9480 2650 9489
rect 2136 9104 2188 9110
rect 2240 9081 2268 9454
rect 2594 9415 2650 9424
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2376 9276 2684 9285
rect 2376 9274 2382 9276
rect 2438 9274 2462 9276
rect 2518 9274 2542 9276
rect 2598 9274 2622 9276
rect 2678 9274 2684 9276
rect 2438 9222 2440 9274
rect 2620 9222 2622 9274
rect 2376 9220 2382 9222
rect 2438 9220 2462 9222
rect 2518 9220 2542 9222
rect 2598 9220 2622 9222
rect 2678 9220 2684 9222
rect 2376 9211 2684 9220
rect 2792 9110 2820 9318
rect 2412 9104 2464 9110
rect 2136 9046 2188 9052
rect 2226 9072 2282 9081
rect 2412 9046 2464 9052
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2226 9007 2282 9016
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8634 2176 8910
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2056 7886 2084 8026
rect 2148 7886 2176 8434
rect 2240 8430 2268 8774
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2332 8276 2360 8774
rect 2424 8566 2452 9046
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2412 8560 2464 8566
rect 2608 8537 2636 8910
rect 2412 8502 2464 8508
rect 2594 8528 2650 8537
rect 2594 8463 2650 8472
rect 2884 8294 2912 9590
rect 3436 9586 3464 9862
rect 3146 9551 3148 9560
rect 3200 9551 3202 9560
rect 3424 9580 3476 9586
rect 3148 9522 3200 9528
rect 3424 9522 3476 9528
rect 3056 9512 3108 9518
rect 2976 9472 3056 9500
rect 2976 9042 3004 9472
rect 3056 9454 3108 9460
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 2976 8480 3004 8978
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3036 8732 3344 8741
rect 3036 8730 3042 8732
rect 3098 8730 3122 8732
rect 3178 8730 3202 8732
rect 3258 8730 3282 8732
rect 3338 8730 3344 8732
rect 3098 8678 3100 8730
rect 3280 8678 3282 8730
rect 3036 8676 3042 8678
rect 3098 8676 3122 8678
rect 3178 8676 3202 8678
rect 3258 8676 3282 8678
rect 3338 8676 3344 8678
rect 3036 8667 3344 8676
rect 3436 8634 3464 8910
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3148 8492 3200 8498
rect 2976 8452 3148 8480
rect 3148 8434 3200 8440
rect 3160 8401 3188 8434
rect 3146 8392 3202 8401
rect 3146 8327 3202 8336
rect 2240 8248 2360 8276
rect 2872 8288 2924 8294
rect 2240 8090 2268 8248
rect 2872 8230 2924 8236
rect 2376 8188 2684 8197
rect 2376 8186 2382 8188
rect 2438 8186 2462 8188
rect 2518 8186 2542 8188
rect 2598 8186 2622 8188
rect 2678 8186 2684 8188
rect 2438 8134 2440 8186
rect 2620 8134 2622 8186
rect 2376 8132 2382 8134
rect 2438 8132 2462 8134
rect 2518 8132 2542 8134
rect 2598 8132 2622 8134
rect 2678 8132 2684 8134
rect 2376 8123 2684 8132
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2884 8022 2912 8230
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 2872 8016 2924 8022
rect 2872 7958 2924 7964
rect 2516 7886 2544 7958
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 3344 7834 3372 8570
rect 3528 8498 3556 9046
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3528 8090 3556 8434
rect 3620 8294 3648 8910
rect 3712 8294 3740 9386
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3804 8634 3832 8910
rect 3792 8628 3844 8634
rect 3792 8570 3844 8576
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3516 8084 3568 8090
rect 3516 8026 3568 8032
rect 2148 7698 2176 7822
rect 2056 7670 2176 7698
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1952 7404 2004 7410
rect 1952 7346 2004 7352
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 6905 1532 7142
rect 1688 7002 1716 7346
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1490 6896 1546 6905
rect 1490 6831 1546 6840
rect 848 6316 900 6322
rect 848 6258 900 6264
rect 860 6089 888 6258
rect 846 6080 902 6089
rect 846 6015 902 6024
rect 1492 5636 1544 5642
rect 1492 5578 1544 5584
rect 1504 5545 1532 5578
rect 1490 5536 1546 5545
rect 1490 5471 1546 5480
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5001 888 5170
rect 2056 5166 2084 7670
rect 2700 7342 2728 7822
rect 3344 7806 3464 7834
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7478 2912 7686
rect 3036 7644 3344 7653
rect 3036 7642 3042 7644
rect 3098 7642 3122 7644
rect 3178 7642 3202 7644
rect 3258 7642 3282 7644
rect 3338 7642 3344 7644
rect 3098 7590 3100 7642
rect 3280 7590 3282 7642
rect 3036 7588 3042 7590
rect 3098 7588 3122 7590
rect 3178 7588 3202 7590
rect 3258 7588 3282 7590
rect 3338 7588 3344 7590
rect 3036 7579 3344 7588
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 2148 6730 2176 7210
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 2240 6662 2268 7142
rect 2376 7100 2684 7109
rect 2376 7098 2382 7100
rect 2438 7098 2462 7100
rect 2518 7098 2542 7100
rect 2598 7098 2622 7100
rect 2678 7098 2684 7100
rect 2438 7046 2440 7098
rect 2620 7046 2622 7098
rect 2376 7044 2382 7046
rect 2438 7044 2462 7046
rect 2518 7044 2542 7046
rect 2598 7044 2622 7046
rect 2678 7044 2684 7046
rect 2376 7035 2684 7044
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2608 6458 2636 6734
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2792 6322 2820 7142
rect 2884 6866 2912 7414
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 2872 6860 2924 6866
rect 2872 6802 2924 6808
rect 3344 6798 3372 7346
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2976 6390 3004 6598
rect 3036 6556 3344 6565
rect 3036 6554 3042 6556
rect 3098 6554 3122 6556
rect 3178 6554 3202 6556
rect 3258 6554 3282 6556
rect 3338 6554 3344 6556
rect 3098 6502 3100 6554
rect 3280 6502 3282 6554
rect 3036 6500 3042 6502
rect 3098 6500 3122 6502
rect 3178 6500 3202 6502
rect 3258 6500 3282 6502
rect 3338 6500 3344 6502
rect 3036 6491 3344 6500
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2376 6012 2684 6021
rect 2376 6010 2382 6012
rect 2438 6010 2462 6012
rect 2518 6010 2542 6012
rect 2598 6010 2622 6012
rect 2678 6010 2684 6012
rect 2438 5958 2440 6010
rect 2620 5958 2622 6010
rect 2376 5956 2382 5958
rect 2438 5956 2462 5958
rect 2518 5956 2542 5958
rect 2598 5956 2622 5958
rect 2678 5956 2684 5958
rect 2376 5947 2684 5956
rect 2688 5704 2740 5710
rect 2792 5692 2820 6054
rect 2884 5710 2912 6190
rect 3160 5914 3188 6190
rect 3436 5914 3464 7806
rect 3712 6730 3740 8230
rect 3804 7410 3832 8434
rect 3896 7886 3924 11154
rect 3988 11150 4016 11290
rect 4080 11218 4108 11698
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4356 11286 4384 11494
rect 4540 11354 4568 12135
rect 4632 11898 4660 13126
rect 5888 13084 6196 13093
rect 5888 13082 5894 13084
rect 5950 13082 5974 13084
rect 6030 13082 6054 13084
rect 6110 13082 6134 13084
rect 6190 13082 6196 13084
rect 5950 13030 5952 13082
rect 6132 13030 6134 13082
rect 5888 13028 5894 13030
rect 5950 13028 5974 13030
rect 6030 13028 6054 13030
rect 6110 13028 6134 13030
rect 6190 13028 6196 13030
rect 5888 13019 6196 13028
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4724 12442 4752 12786
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 12442 4844 12718
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 5000 12306 5028 12786
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5228 12540 5536 12549
rect 5228 12538 5234 12540
rect 5290 12538 5314 12540
rect 5370 12538 5394 12540
rect 5450 12538 5474 12540
rect 5530 12538 5536 12540
rect 5290 12486 5292 12538
rect 5472 12486 5474 12538
rect 5228 12484 5234 12486
rect 5290 12484 5314 12486
rect 5370 12484 5394 12486
rect 5450 12484 5474 12486
rect 5530 12484 5536 12486
rect 5228 12475 5536 12484
rect 5828 12374 5856 12718
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 5172 12300 5224 12306
rect 5172 12242 5224 12248
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4528 11348 4580 11354
rect 4528 11290 4580 11296
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4080 10606 4108 11018
rect 4172 10674 4200 11018
rect 4356 10810 4384 11222
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 8634 4016 9454
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 3988 8430 4016 8570
rect 4080 8498 4108 10542
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4172 9722 4200 10406
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4264 9081 4292 9114
rect 4250 9072 4306 9081
rect 4160 9036 4212 9042
rect 4250 9007 4306 9016
rect 4160 8978 4212 8984
rect 4172 8634 4200 8978
rect 4540 8974 4568 11290
rect 4632 11234 4660 11834
rect 4816 11558 4844 12174
rect 5080 12164 5132 12170
rect 5080 12106 5132 12112
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4632 11206 4752 11234
rect 4632 10674 4660 11206
rect 4724 11150 4752 11206
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 4908 11082 4936 11834
rect 5092 11354 5120 12106
rect 5184 11898 5212 12242
rect 5262 12200 5318 12209
rect 5262 12135 5318 12144
rect 5540 12164 5592 12170
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5276 11830 5304 12135
rect 5540 12106 5592 12112
rect 5264 11824 5316 11830
rect 5264 11766 5316 11772
rect 5552 11762 5580 12106
rect 5888 11996 6196 12005
rect 5888 11994 5894 11996
rect 5950 11994 5974 11996
rect 6030 11994 6054 11996
rect 6110 11994 6134 11996
rect 6190 11994 6196 11996
rect 5950 11942 5952 11994
rect 6132 11942 6134 11994
rect 5888 11940 5894 11942
rect 5950 11940 5974 11942
rect 6030 11940 6054 11942
rect 6110 11940 6134 11942
rect 6190 11940 6196 11942
rect 5888 11931 6196 11940
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5228 11452 5536 11461
rect 5228 11450 5234 11452
rect 5290 11450 5314 11452
rect 5370 11450 5394 11452
rect 5450 11450 5474 11452
rect 5530 11450 5536 11452
rect 5290 11398 5292 11450
rect 5472 11398 5474 11450
rect 5228 11396 5234 11398
rect 5290 11396 5314 11398
rect 5370 11396 5394 11398
rect 5450 11396 5474 11398
rect 5530 11396 5536 11398
rect 5228 11387 5536 11396
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5644 11082 5672 11494
rect 5736 11354 5764 11630
rect 6288 11626 6316 13126
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6748 12306 6776 12582
rect 7116 12442 7144 12786
rect 7104 12436 7156 12442
rect 7104 12378 7156 12384
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6840 12170 6868 12310
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 6288 11082 6316 11562
rect 6656 11286 6684 11698
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6840 11082 6868 12106
rect 7012 11348 7064 11354
rect 7208 11336 7236 13126
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7668 12442 7696 12786
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7668 11898 7696 12378
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7852 11762 7880 13194
rect 8740 13084 9048 13093
rect 8740 13082 8746 13084
rect 8802 13082 8826 13084
rect 8882 13082 8906 13084
rect 8962 13082 8986 13084
rect 9042 13082 9048 13084
rect 8802 13030 8804 13082
rect 8984 13030 8986 13082
rect 8740 13028 8746 13030
rect 8802 13028 8826 13030
rect 8882 13028 8906 13030
rect 8962 13028 8986 13030
rect 9042 13028 9048 13030
rect 8740 13019 9048 13028
rect 11592 13084 11900 13093
rect 11592 13082 11598 13084
rect 11654 13082 11678 13084
rect 11734 13082 11758 13084
rect 11814 13082 11838 13084
rect 11894 13082 11900 13084
rect 11654 13030 11656 13082
rect 11836 13030 11838 13082
rect 11592 13028 11598 13030
rect 11654 13028 11678 13030
rect 11734 13028 11758 13030
rect 11814 13028 11838 13030
rect 11894 13028 11900 13030
rect 11592 13019 11900 13028
rect 9036 12844 9088 12850
rect 9036 12786 9088 12792
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 7944 12238 7972 12718
rect 8080 12540 8388 12549
rect 8080 12538 8086 12540
rect 8142 12538 8166 12540
rect 8222 12538 8246 12540
rect 8302 12538 8326 12540
rect 8382 12538 8388 12540
rect 8142 12486 8144 12538
rect 8324 12486 8326 12538
rect 8080 12484 8086 12486
rect 8142 12484 8166 12486
rect 8222 12484 8246 12486
rect 8302 12484 8326 12486
rect 8382 12484 8388 12486
rect 8080 12475 8388 12484
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 7932 12232 7984 12238
rect 7932 12174 7984 12180
rect 8680 11898 8708 12378
rect 8956 12238 8984 12718
rect 9048 12442 9076 12786
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 8740 11996 9048 12005
rect 8740 11994 8746 11996
rect 8802 11994 8826 11996
rect 8882 11994 8906 11996
rect 8962 11994 8986 11996
rect 9042 11994 9048 11996
rect 8802 11942 8804 11994
rect 8984 11942 8986 11994
rect 8740 11940 8746 11942
rect 8802 11940 8826 11942
rect 8882 11940 8906 11942
rect 8962 11940 8986 11942
rect 9042 11940 9048 11942
rect 8740 11931 9048 11940
rect 9324 11898 9352 12038
rect 9600 11898 9628 12038
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9692 11778 9720 12378
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 9600 11762 9720 11778
rect 9968 11762 9996 12038
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 9588 11756 9720 11762
rect 9640 11750 9720 11756
rect 9956 11756 10008 11762
rect 9588 11698 9640 11704
rect 9956 11698 10008 11704
rect 7300 11558 7328 11698
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7064 11308 7236 11336
rect 7012 11290 7064 11296
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 4908 10810 4936 11018
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4724 9432 4752 10202
rect 4816 9654 4844 10474
rect 5092 10470 5120 10950
rect 5644 10810 5672 11018
rect 5888 10908 6196 10917
rect 5888 10906 5894 10908
rect 5950 10906 5974 10908
rect 6030 10906 6054 10908
rect 6110 10906 6134 10908
rect 6190 10906 6196 10908
rect 5950 10854 5952 10906
rect 6132 10854 6134 10906
rect 5888 10852 5894 10854
rect 5950 10852 5974 10854
rect 6030 10852 6054 10854
rect 6110 10852 6134 10854
rect 6190 10852 6196 10854
rect 5888 10843 6196 10852
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 6288 10742 6316 11018
rect 6276 10736 6328 10742
rect 6276 10678 6328 10684
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4804 9648 4856 9654
rect 4804 9590 4856 9596
rect 4804 9444 4856 9450
rect 4724 9404 4804 9432
rect 4804 9386 4856 9392
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 3884 7880 3936 7886
rect 3884 7822 3936 7828
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3896 7274 3924 7822
rect 3988 7818 4016 8366
rect 4448 8090 4476 8434
rect 4540 8401 4568 8910
rect 4526 8392 4582 8401
rect 4526 8327 4528 8336
rect 4580 8327 4582 8336
rect 4528 8298 4580 8304
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4540 7886 4568 8298
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 3976 7812 4028 7818
rect 3976 7754 4028 7760
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3700 6724 3752 6730
rect 3700 6666 3752 6672
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 2740 5664 2820 5692
rect 2688 5646 2740 5652
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 2240 5302 2268 5578
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 846 4992 902 5001
rect 846 4927 902 4936
rect 2240 4622 2268 5238
rect 2792 5234 2820 5664
rect 2872 5704 2924 5710
rect 2872 5646 2924 5652
rect 2884 5574 2912 5646
rect 3436 5574 3464 5850
rect 3712 5846 3740 6666
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6186 3832 6598
rect 3792 6180 3844 6186
rect 3792 6122 3844 6128
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2376 4924 2684 4933
rect 2376 4922 2382 4924
rect 2438 4922 2462 4924
rect 2518 4922 2542 4924
rect 2598 4922 2622 4924
rect 2678 4922 2684 4924
rect 2438 4870 2440 4922
rect 2620 4870 2622 4922
rect 2376 4868 2382 4870
rect 2438 4868 2462 4870
rect 2518 4868 2542 4870
rect 2598 4868 2622 4870
rect 2678 4868 2684 4870
rect 2376 4859 2684 4868
rect 2884 4826 2912 5510
rect 3036 5468 3344 5477
rect 3036 5466 3042 5468
rect 3098 5466 3122 5468
rect 3178 5466 3202 5468
rect 3258 5466 3282 5468
rect 3338 5466 3344 5468
rect 3098 5414 3100 5466
rect 3280 5414 3282 5466
rect 3036 5412 3042 5414
rect 3098 5412 3122 5414
rect 3178 5412 3202 5414
rect 3258 5412 3282 5414
rect 3338 5412 3344 5414
rect 3036 5403 3344 5412
rect 3528 5234 3556 5714
rect 3988 5710 4016 7414
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4080 5710 4108 6258
rect 4724 5914 4752 6258
rect 4816 6118 4844 9386
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4894 8528 4950 8537
rect 4894 8463 4896 8472
rect 4948 8463 4950 8472
rect 4896 8434 4948 8440
rect 4908 6798 4936 8434
rect 5000 7954 5028 9046
rect 5092 8548 5120 10406
rect 5228 10364 5536 10373
rect 5228 10362 5234 10364
rect 5290 10362 5314 10364
rect 5370 10362 5394 10364
rect 5450 10362 5474 10364
rect 5530 10362 5536 10364
rect 5290 10310 5292 10362
rect 5472 10310 5474 10362
rect 5228 10308 5234 10310
rect 5290 10308 5314 10310
rect 5370 10308 5394 10310
rect 5450 10308 5474 10310
rect 5530 10308 5536 10310
rect 5228 10299 5536 10308
rect 6840 10062 6868 11018
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10470 6960 10950
rect 7024 10674 7052 11290
rect 7576 11218 7604 11630
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7208 10810 7236 11154
rect 7656 11144 7708 11150
rect 7654 11112 7656 11121
rect 7760 11132 7788 11494
rect 7852 11234 7880 11698
rect 8484 11688 8536 11694
rect 8484 11630 8536 11636
rect 8080 11452 8388 11461
rect 8080 11450 8086 11452
rect 8142 11450 8166 11452
rect 8222 11450 8246 11452
rect 8302 11450 8326 11452
rect 8382 11450 8388 11452
rect 8142 11398 8144 11450
rect 8324 11398 8326 11450
rect 8080 11396 8086 11398
rect 8142 11396 8166 11398
rect 8222 11396 8246 11398
rect 8302 11396 8326 11398
rect 8382 11396 8388 11398
rect 8080 11387 8388 11396
rect 8496 11354 8524 11630
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 7852 11206 7972 11234
rect 7944 11150 7972 11206
rect 7840 11144 7892 11150
rect 7708 11112 7710 11121
rect 7760 11104 7840 11132
rect 7840 11086 7892 11092
rect 7932 11144 7984 11150
rect 8484 11144 8536 11150
rect 7932 11086 7984 11092
rect 8482 11112 8484 11121
rect 8536 11112 8538 11121
rect 7654 11047 7710 11056
rect 7380 11008 7432 11014
rect 7380 10950 7432 10956
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 5888 9820 6196 9829
rect 5888 9818 5894 9820
rect 5950 9818 5974 9820
rect 6030 9818 6054 9820
rect 6110 9818 6134 9820
rect 6190 9818 6196 9820
rect 5950 9766 5952 9818
rect 6132 9766 6134 9818
rect 5888 9764 5894 9766
rect 5950 9764 5974 9766
rect 6030 9764 6054 9766
rect 6110 9764 6134 9766
rect 6190 9764 6196 9766
rect 5888 9755 6196 9764
rect 6840 9722 6868 9998
rect 6932 9926 6960 10406
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5228 9276 5536 9285
rect 5228 9274 5234 9276
rect 5290 9274 5314 9276
rect 5370 9274 5394 9276
rect 5450 9274 5474 9276
rect 5530 9274 5536 9276
rect 5290 9222 5292 9274
rect 5472 9222 5474 9274
rect 5228 9220 5234 9222
rect 5290 9220 5314 9222
rect 5370 9220 5394 9222
rect 5450 9220 5474 9222
rect 5530 9220 5536 9222
rect 5228 9211 5536 9220
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5276 8566 5304 8910
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5264 8560 5316 8566
rect 5092 8520 5264 8548
rect 4988 7948 5040 7954
rect 4988 7890 5040 7896
rect 5092 7886 5120 8520
rect 5264 8502 5316 8508
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5368 8294 5396 8434
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5228 8188 5536 8197
rect 5228 8186 5234 8188
rect 5290 8186 5314 8188
rect 5370 8186 5394 8188
rect 5450 8186 5474 8188
rect 5530 8186 5536 8188
rect 5290 8134 5292 8186
rect 5472 8134 5474 8186
rect 5228 8132 5234 8134
rect 5290 8132 5314 8134
rect 5370 8132 5394 8134
rect 5450 8132 5474 8134
rect 5530 8132 5536 8134
rect 5228 8123 5536 8132
rect 5644 7886 5672 8570
rect 5736 8294 5764 9522
rect 6932 9518 6960 9862
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 6092 9376 6144 9382
rect 6092 9318 6144 9324
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 5828 9178 5856 9318
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5920 8820 5948 9318
rect 6104 9110 6132 9318
rect 6092 9104 6144 9110
rect 6092 9046 6144 9052
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 5828 8792 5948 8820
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6458 4936 6734
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4724 5710 4752 5850
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 4068 5704 4120 5710
rect 4436 5704 4488 5710
rect 4068 5646 4120 5652
rect 4158 5672 4214 5681
rect 4080 5370 4108 5646
rect 4436 5646 4488 5652
rect 4712 5704 4764 5710
rect 4712 5646 4764 5652
rect 4896 5704 4948 5710
rect 5000 5692 5028 6190
rect 4948 5664 5028 5692
rect 4896 5646 4948 5652
rect 4158 5607 4160 5616
rect 4212 5607 4214 5616
rect 4160 5578 4212 5584
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3252 4826 3280 5170
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3528 4622 3556 5170
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3036 4380 3344 4389
rect 3036 4378 3042 4380
rect 3098 4378 3122 4380
rect 3178 4378 3202 4380
rect 3258 4378 3282 4380
rect 3338 4378 3344 4380
rect 3098 4326 3100 4378
rect 3280 4326 3282 4378
rect 3036 4324 3042 4326
rect 3098 4324 3122 4326
rect 3178 4324 3202 4326
rect 3258 4324 3282 4326
rect 3338 4324 3344 4326
rect 3036 4315 3344 4324
rect 4080 4214 4108 4762
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4172 3942 4200 4558
rect 4356 4146 4384 5510
rect 4448 5302 4476 5646
rect 4528 5636 4580 5642
rect 4528 5578 4580 5584
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 4448 4690 4476 5238
rect 4436 4684 4488 4690
rect 4436 4626 4488 4632
rect 4448 4282 4476 4626
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 4160 3936 4212 3942
rect 4160 3878 4212 3884
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 2376 3836 2684 3845
rect 2376 3834 2382 3836
rect 2438 3834 2462 3836
rect 2518 3834 2542 3836
rect 2598 3834 2622 3836
rect 2678 3834 2684 3836
rect 2438 3782 2440 3834
rect 2620 3782 2622 3834
rect 2376 3780 2382 3782
rect 2438 3780 2462 3782
rect 2518 3780 2542 3782
rect 2598 3780 2622 3782
rect 2678 3780 2684 3782
rect 2376 3771 2684 3780
rect 4356 3618 4384 3878
rect 4448 3738 4476 4014
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4356 3590 4476 3618
rect 4448 3534 4476 3590
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4344 3528 4396 3534
rect 4344 3470 4396 3476
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 3036 3292 3344 3301
rect 3036 3290 3042 3292
rect 3098 3290 3122 3292
rect 3178 3290 3202 3292
rect 3258 3290 3282 3292
rect 3338 3290 3344 3292
rect 3098 3238 3100 3290
rect 3280 3238 3282 3290
rect 3036 3236 3042 3238
rect 3098 3236 3122 3238
rect 3178 3236 3202 3238
rect 3258 3236 3282 3238
rect 3338 3236 3344 3238
rect 3036 3227 3344 3236
rect 4172 3058 4200 3470
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4356 2990 4384 3470
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 2376 2748 2684 2757
rect 2376 2746 2382 2748
rect 2438 2746 2462 2748
rect 2518 2746 2542 2748
rect 2598 2746 2622 2748
rect 2678 2746 2684 2748
rect 2438 2694 2440 2746
rect 2620 2694 2622 2746
rect 2376 2692 2382 2694
rect 2438 2692 2462 2694
rect 2518 2692 2542 2694
rect 2598 2692 2622 2694
rect 2678 2692 2684 2694
rect 2376 2683 2684 2692
rect 4540 2446 4568 5578
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 2446 4660 3878
rect 4724 3058 4752 5646
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4816 4826 4844 5170
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 5000 4622 5028 5664
rect 5092 5522 5120 7686
rect 5228 7100 5536 7109
rect 5228 7098 5234 7100
rect 5290 7098 5314 7100
rect 5370 7098 5394 7100
rect 5450 7098 5474 7100
rect 5530 7098 5536 7100
rect 5290 7046 5292 7098
rect 5472 7046 5474 7098
rect 5228 7044 5234 7046
rect 5290 7044 5314 7046
rect 5370 7044 5394 7046
rect 5450 7044 5474 7046
rect 5530 7044 5536 7046
rect 5228 7035 5536 7044
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5368 6662 5396 6870
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5184 6322 5212 6598
rect 5828 6322 5856 8792
rect 5888 8732 6196 8741
rect 5888 8730 5894 8732
rect 5950 8730 5974 8732
rect 6030 8730 6054 8732
rect 6110 8730 6134 8732
rect 6190 8730 6196 8732
rect 5950 8678 5952 8730
rect 6132 8678 6134 8730
rect 5888 8676 5894 8678
rect 5950 8676 5974 8678
rect 6030 8676 6054 8678
rect 6110 8676 6134 8678
rect 6190 8676 6196 8678
rect 5888 8667 6196 8676
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5920 8090 5948 8434
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5888 7644 6196 7653
rect 5888 7642 5894 7644
rect 5950 7642 5974 7644
rect 6030 7642 6054 7644
rect 6110 7642 6134 7644
rect 6190 7642 6196 7644
rect 5950 7590 5952 7642
rect 6132 7590 6134 7642
rect 5888 7588 5894 7590
rect 5950 7588 5974 7590
rect 6030 7588 6054 7590
rect 6110 7588 6134 7590
rect 6190 7588 6196 7590
rect 5888 7579 6196 7588
rect 6288 6662 6316 8978
rect 6748 8974 6776 9318
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6840 8430 6868 9318
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 5888 6556 6196 6565
rect 5888 6554 5894 6556
rect 5950 6554 5974 6556
rect 6030 6554 6054 6556
rect 6110 6554 6134 6556
rect 6190 6554 6196 6556
rect 5950 6502 5952 6554
rect 6132 6502 6134 6554
rect 5888 6500 5894 6502
rect 5950 6500 5974 6502
rect 6030 6500 6054 6502
rect 6110 6500 6134 6502
rect 6190 6500 6196 6502
rect 5888 6491 6196 6500
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5460 6186 5764 6202
rect 5448 6180 5764 6186
rect 5500 6174 5764 6180
rect 5448 6122 5500 6128
rect 5632 6112 5684 6118
rect 5632 6054 5684 6060
rect 5228 6012 5536 6021
rect 5228 6010 5234 6012
rect 5290 6010 5314 6012
rect 5370 6010 5394 6012
rect 5450 6010 5474 6012
rect 5530 6010 5536 6012
rect 5290 5958 5292 6010
rect 5472 5958 5474 6010
rect 5228 5956 5234 5958
rect 5290 5956 5314 5958
rect 5370 5956 5394 5958
rect 5450 5956 5474 5958
rect 5530 5956 5536 5958
rect 5228 5947 5536 5956
rect 5644 5914 5672 6054
rect 5736 5914 5764 6174
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 6012 5710 6040 5850
rect 5816 5704 5868 5710
rect 6000 5704 6052 5710
rect 5816 5646 5868 5652
rect 5998 5672 6000 5681
rect 6052 5672 6054 5681
rect 5172 5568 5224 5574
rect 5092 5516 5172 5522
rect 5092 5510 5224 5516
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5092 5494 5212 5510
rect 5092 5302 5120 5494
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 5228 4924 5536 4933
rect 5228 4922 5234 4924
rect 5290 4922 5314 4924
rect 5370 4922 5394 4924
rect 5450 4922 5474 4924
rect 5530 4922 5536 4924
rect 5290 4870 5292 4922
rect 5472 4870 5474 4922
rect 5228 4868 5234 4870
rect 5290 4868 5314 4870
rect 5370 4868 5394 4870
rect 5450 4868 5474 4870
rect 5530 4868 5536 4870
rect 5228 4859 5536 4868
rect 5644 4808 5672 5510
rect 5552 4780 5672 4808
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5000 4214 5028 4558
rect 4988 4208 5040 4214
rect 4988 4150 5040 4156
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4816 3738 4844 4014
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 5000 2650 5028 4150
rect 5092 4078 5120 4558
rect 5552 4282 5580 4780
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 5092 3194 5120 4014
rect 5228 3836 5536 3845
rect 5228 3834 5234 3836
rect 5290 3834 5314 3836
rect 5370 3834 5394 3836
rect 5450 3834 5474 3836
rect 5530 3834 5536 3836
rect 5290 3782 5292 3834
rect 5472 3782 5474 3834
rect 5228 3780 5234 3782
rect 5290 3780 5314 3782
rect 5370 3780 5394 3782
rect 5450 3780 5474 3782
rect 5530 3780 5536 3782
rect 5228 3771 5536 3780
rect 5644 3670 5672 4422
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5632 3664 5684 3670
rect 5632 3606 5684 3612
rect 5356 3528 5408 3534
rect 5644 3516 5672 3606
rect 5736 3602 5764 4150
rect 5828 4010 5856 5646
rect 5998 5607 6054 5616
rect 6288 5574 6316 6598
rect 6380 6390 6408 8298
rect 6552 7948 6604 7954
rect 6552 7890 6604 7896
rect 6564 7546 6592 7890
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6748 7410 6776 7822
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6380 5914 6408 6326
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 5888 5468 6196 5477
rect 5888 5466 5894 5468
rect 5950 5466 5974 5468
rect 6030 5466 6054 5468
rect 6110 5466 6134 5468
rect 6190 5466 6196 5468
rect 5950 5414 5952 5466
rect 6132 5414 6134 5466
rect 5888 5412 5894 5414
rect 5950 5412 5974 5414
rect 6030 5412 6054 5414
rect 6110 5412 6134 5414
rect 6190 5412 6196 5414
rect 5888 5403 6196 5412
rect 6380 4622 6408 5850
rect 6564 5166 6592 7346
rect 7024 7342 7052 10610
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7116 9586 7144 10134
rect 7208 9722 7236 10746
rect 7392 10062 7420 10950
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7208 9058 7236 9658
rect 7392 9654 7420 9998
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7668 9586 7696 9862
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7116 9030 7236 9058
rect 7564 9036 7616 9042
rect 7116 8634 7144 9030
rect 7564 8978 7616 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7116 7886 7144 8570
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7024 6934 7052 7278
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 7208 6730 7236 8230
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7116 6322 7144 6394
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7116 5710 7144 6258
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 5888 4380 6196 4389
rect 5888 4378 5894 4380
rect 5950 4378 5974 4380
rect 6030 4378 6054 4380
rect 6110 4378 6134 4380
rect 6190 4378 6196 4380
rect 5950 4326 5952 4378
rect 6132 4326 6134 4378
rect 5888 4324 5894 4326
rect 5950 4324 5974 4326
rect 6030 4324 6054 4326
rect 6110 4324 6134 4326
rect 6190 4324 6196 4326
rect 5888 4315 6196 4324
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6012 3738 6040 3878
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5408 3488 5672 3516
rect 5356 3470 5408 3476
rect 5736 3466 5764 3538
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 5736 3194 5764 3402
rect 5828 3194 5856 3402
rect 5888 3292 6196 3301
rect 5888 3290 5894 3292
rect 5950 3290 5974 3292
rect 6030 3290 6054 3292
rect 6110 3290 6134 3292
rect 6190 3290 6196 3292
rect 5950 3238 5952 3290
rect 6132 3238 6134 3290
rect 5888 3236 5894 3238
rect 5950 3236 5974 3238
rect 6030 3236 6054 3238
rect 6110 3236 6134 3238
rect 6190 3236 6196 3238
rect 5888 3227 6196 3236
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6288 3058 6316 3402
rect 6380 3058 6408 4014
rect 6460 3664 6512 3670
rect 6460 3606 6512 3612
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 5644 2774 5672 2994
rect 6288 2854 6316 2994
rect 6472 2990 6500 3606
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6564 2922 6592 3334
rect 6840 2922 6868 4082
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6932 2990 6960 3538
rect 7024 3466 7052 4966
rect 7116 4554 7144 5170
rect 7208 5166 7236 6666
rect 7392 6458 7420 8910
rect 7472 7268 7524 7274
rect 7472 7210 7524 7216
rect 7484 7002 7512 7210
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 5710 7420 6190
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7300 5370 7328 5646
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7104 4548 7156 4554
rect 7104 4490 7156 4496
rect 7116 3534 7144 4490
rect 7484 3534 7512 6598
rect 7576 5710 7604 8978
rect 7668 8906 7696 9522
rect 7760 9042 7788 9590
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7656 8900 7708 8906
rect 7656 8842 7708 8848
rect 7760 8362 7788 8978
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7944 7834 7972 11086
rect 8482 11047 8538 11056
rect 8080 10364 8388 10373
rect 8080 10362 8086 10364
rect 8142 10362 8166 10364
rect 8222 10362 8246 10364
rect 8302 10362 8326 10364
rect 8382 10362 8388 10364
rect 8142 10310 8144 10362
rect 8324 10310 8326 10362
rect 8080 10308 8086 10310
rect 8142 10308 8166 10310
rect 8222 10308 8246 10310
rect 8302 10308 8326 10310
rect 8382 10308 8388 10310
rect 8080 10299 8388 10308
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8080 9276 8388 9285
rect 8080 9274 8086 9276
rect 8142 9274 8166 9276
rect 8222 9274 8246 9276
rect 8302 9274 8326 9276
rect 8382 9274 8388 9276
rect 8142 9222 8144 9274
rect 8324 9222 8326 9274
rect 8080 9220 8086 9222
rect 8142 9220 8166 9222
rect 8222 9220 8246 9222
rect 8302 9220 8326 9222
rect 8382 9220 8388 9222
rect 8080 9211 8388 9220
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8036 8634 8064 8910
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8128 8566 8156 8842
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8312 8294 8340 8910
rect 8496 8498 8524 9318
rect 8588 9110 8616 11494
rect 8740 10908 9048 10917
rect 8740 10906 8746 10908
rect 8802 10906 8826 10908
rect 8882 10906 8906 10908
rect 8962 10906 8986 10908
rect 9042 10906 9048 10908
rect 8802 10854 8804 10906
rect 8984 10854 8986 10906
rect 8740 10852 8746 10854
rect 8802 10852 8826 10854
rect 8882 10852 8906 10854
rect 8962 10852 8986 10854
rect 9042 10852 9048 10854
rect 8740 10843 9048 10852
rect 10244 10674 10272 12582
rect 10336 12238 10364 12650
rect 10932 12540 11240 12549
rect 10932 12538 10938 12540
rect 10994 12538 11018 12540
rect 11074 12538 11098 12540
rect 11154 12538 11178 12540
rect 11234 12538 11240 12540
rect 10994 12486 10996 12538
rect 11176 12486 11178 12538
rect 10932 12484 10938 12486
rect 10994 12484 11018 12486
rect 11074 12484 11098 12486
rect 11154 12484 11178 12486
rect 11234 12484 11240 12486
rect 10932 12475 11240 12484
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10612 11150 10640 11494
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10704 10826 10732 11290
rect 10796 11150 10824 12310
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11532 11830 11560 12038
rect 11592 11996 11900 12005
rect 11592 11994 11598 11996
rect 11654 11994 11678 11996
rect 11734 11994 11758 11996
rect 11814 11994 11838 11996
rect 11894 11994 11900 11996
rect 11654 11942 11656 11994
rect 11836 11942 11838 11994
rect 11592 11940 11598 11942
rect 11654 11940 11678 11942
rect 11734 11940 11758 11942
rect 11814 11940 11838 11942
rect 11894 11940 11900 11942
rect 11592 11931 11900 11940
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 10932 11452 11240 11461
rect 10932 11450 10938 11452
rect 10994 11450 11018 11452
rect 11074 11450 11098 11452
rect 11154 11450 11178 11452
rect 11234 11450 11240 11452
rect 10994 11398 10996 11450
rect 11176 11398 11178 11450
rect 10932 11396 10938 11398
rect 10994 11396 11018 11398
rect 11074 11396 11098 11398
rect 11154 11396 11178 11398
rect 11234 11396 11240 11398
rect 10932 11387 11240 11396
rect 11532 11218 11560 11766
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10612 10798 10732 10826
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10244 10266 10272 10610
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 8740 9820 9048 9829
rect 8740 9818 8746 9820
rect 8802 9818 8826 9820
rect 8882 9818 8906 9820
rect 8962 9818 8986 9820
rect 9042 9818 9048 9820
rect 8802 9766 8804 9818
rect 8984 9766 8986 9818
rect 8740 9764 8746 9766
rect 8802 9764 8826 9766
rect 8882 9764 8906 9766
rect 8962 9764 8986 9766
rect 9042 9764 9048 9766
rect 8740 9755 9048 9764
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8080 8188 8388 8197
rect 8080 8186 8086 8188
rect 8142 8186 8166 8188
rect 8222 8186 8246 8188
rect 8302 8186 8326 8188
rect 8382 8186 8388 8188
rect 8142 8134 8144 8186
rect 8324 8134 8326 8186
rect 8080 8132 8086 8134
rect 8142 8132 8166 8134
rect 8222 8132 8246 8134
rect 8302 8132 8326 8134
rect 8382 8132 8388 8134
rect 8080 8123 8388 8132
rect 8116 7880 8168 7886
rect 7944 7806 8064 7834
rect 8116 7822 8168 7828
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7944 7410 7972 7686
rect 8036 7410 8064 7806
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7852 6798 7880 7278
rect 7944 6866 7972 7346
rect 8128 7342 8156 7822
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8080 7100 8388 7109
rect 8080 7098 8086 7100
rect 8142 7098 8166 7100
rect 8222 7098 8246 7100
rect 8302 7098 8326 7100
rect 8382 7098 8388 7100
rect 8142 7046 8144 7098
rect 8324 7046 8326 7098
rect 8080 7044 8086 7046
rect 8142 7044 8166 7046
rect 8222 7044 8246 7046
rect 8302 7044 8326 7046
rect 8382 7044 8388 7046
rect 8080 7035 8388 7044
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 8496 6798 8524 7142
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6322 8524 6598
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8080 6012 8388 6021
rect 8080 6010 8086 6012
rect 8142 6010 8166 6012
rect 8222 6010 8246 6012
rect 8302 6010 8326 6012
rect 8382 6010 8388 6012
rect 8142 5958 8144 6010
rect 8324 5958 8326 6010
rect 8080 5956 8086 5958
rect 8142 5956 8166 5958
rect 8222 5956 8246 5958
rect 8302 5956 8326 5958
rect 8382 5956 8388 5958
rect 8080 5947 8388 5956
rect 8588 5710 8616 6190
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8680 5642 8708 9522
rect 9770 9480 9826 9489
rect 9128 9444 9180 9450
rect 9770 9415 9826 9424
rect 9128 9386 9180 9392
rect 9140 8974 9168 9386
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9416 8922 9444 8978
rect 9784 8974 9812 9415
rect 10244 9178 10272 9998
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10324 9104 10376 9110
rect 10244 9052 10324 9058
rect 10244 9046 10376 9052
rect 10244 9030 10364 9046
rect 9772 8968 9824 8974
rect 8740 8732 9048 8741
rect 8740 8730 8746 8732
rect 8802 8730 8826 8732
rect 8882 8730 8906 8732
rect 8962 8730 8986 8732
rect 9042 8730 9048 8732
rect 8802 8678 8804 8730
rect 8984 8678 8986 8730
rect 8740 8676 8746 8678
rect 8802 8676 8826 8678
rect 8882 8676 8906 8678
rect 8962 8676 8986 8678
rect 9042 8676 9048 8678
rect 8740 8667 9048 8676
rect 9140 8498 9168 8910
rect 9416 8894 9536 8922
rect 9772 8910 9824 8916
rect 9508 8498 9536 8894
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9600 8634 9628 8774
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9784 8498 9812 8774
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9508 8090 9536 8434
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9496 8084 9548 8090
rect 9496 8026 9548 8032
rect 8740 7644 9048 7653
rect 8740 7642 8746 7644
rect 8802 7642 8826 7644
rect 8882 7642 8906 7644
rect 8962 7642 8986 7644
rect 9042 7642 9048 7644
rect 8802 7590 8804 7642
rect 8984 7590 8986 7642
rect 8740 7588 8746 7590
rect 8802 7588 8826 7590
rect 8882 7588 8906 7590
rect 8962 7588 8986 7590
rect 9042 7588 9048 7590
rect 8740 7579 9048 7588
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 8740 6556 9048 6565
rect 8740 6554 8746 6556
rect 8802 6554 8826 6556
rect 8882 6554 8906 6556
rect 8962 6554 8986 6556
rect 9042 6554 9048 6556
rect 8802 6502 8804 6554
rect 8984 6502 8986 6554
rect 8740 6500 8746 6502
rect 8802 6500 8826 6502
rect 8882 6500 8906 6502
rect 8962 6500 8986 6502
rect 9042 6500 9048 6502
rect 8740 6491 9048 6500
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 9048 5914 9076 6258
rect 9232 6186 9260 6666
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6390 9536 6598
rect 9496 6384 9548 6390
rect 9496 6326 9548 6332
rect 9876 6225 9904 8366
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9968 6798 9996 7142
rect 10048 6928 10100 6934
rect 10048 6870 10100 6876
rect 10060 6798 10088 6870
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9862 6216 9918 6225
rect 9220 6180 9272 6186
rect 9862 6151 9918 6160
rect 9220 6122 9272 6128
rect 9036 5908 9088 5914
rect 9036 5850 9088 5856
rect 9232 5778 9260 6122
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5778 9812 6054
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7668 4826 7696 5102
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7760 4146 7788 5510
rect 8576 5296 8628 5302
rect 8680 5250 8708 5578
rect 8740 5468 9048 5477
rect 8740 5466 8746 5468
rect 8802 5466 8826 5468
rect 8882 5466 8906 5468
rect 8962 5466 8986 5468
rect 9042 5466 9048 5468
rect 8802 5414 8804 5466
rect 8984 5414 8986 5466
rect 8740 5412 8746 5414
rect 8802 5412 8826 5414
rect 8882 5412 8906 5414
rect 8962 5412 8986 5414
rect 9042 5412 9048 5414
rect 8740 5403 9048 5412
rect 8628 5244 8708 5250
rect 8576 5238 8708 5244
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8588 5222 8708 5238
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7852 4826 7880 5102
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7944 4622 7972 5170
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8080 4924 8388 4933
rect 8080 4922 8086 4924
rect 8142 4922 8166 4924
rect 8222 4922 8246 4924
rect 8302 4922 8326 4924
rect 8382 4922 8388 4924
rect 8142 4870 8144 4922
rect 8324 4870 8326 4922
rect 8080 4868 8086 4870
rect 8142 4868 8166 4870
rect 8222 4868 8246 4870
rect 8302 4868 8326 4870
rect 8382 4868 8388 4870
rect 8080 4859 8388 4868
rect 8496 4826 8524 5102
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8588 4706 8616 5222
rect 8312 4678 8616 4706
rect 8312 4622 8340 4678
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7944 4146 7972 4558
rect 8588 4554 8616 4678
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8740 4380 9048 4389
rect 8740 4378 8746 4380
rect 8802 4378 8826 4380
rect 8882 4378 8906 4380
rect 8962 4378 8986 4380
rect 9042 4378 9048 4380
rect 8802 4326 8804 4378
rect 8984 4326 8986 4378
rect 8740 4324 8746 4326
rect 8802 4324 8826 4326
rect 8882 4324 8906 4326
rect 8962 4324 8986 4326
rect 9042 4324 9048 4326
rect 8740 4315 9048 4324
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 7116 3346 7144 3470
rect 7024 3318 7144 3346
rect 7024 3058 7052 3318
rect 7576 3194 7604 4014
rect 7564 3188 7616 3194
rect 7564 3130 7616 3136
rect 7944 3058 7972 4082
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 8080 3836 8388 3845
rect 8080 3834 8086 3836
rect 8142 3834 8166 3836
rect 8222 3834 8246 3836
rect 8302 3834 8326 3836
rect 8382 3834 8388 3836
rect 8142 3782 8144 3834
rect 8324 3782 8326 3834
rect 8080 3780 8086 3782
rect 8142 3780 8166 3782
rect 8222 3780 8246 3782
rect 8302 3780 8326 3782
rect 8382 3780 8388 3782
rect 8080 3771 8388 3780
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 6920 2984 6972 2990
rect 6920 2926 6972 2932
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6828 2916 6880 2922
rect 6828 2858 6880 2864
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 5228 2748 5536 2757
rect 5228 2746 5234 2748
rect 5290 2746 5314 2748
rect 5370 2746 5394 2748
rect 5450 2746 5474 2748
rect 5530 2746 5536 2748
rect 5644 2746 5764 2774
rect 5290 2694 5292 2746
rect 5472 2694 5474 2746
rect 5228 2692 5234 2694
rect 5290 2692 5314 2694
rect 5370 2692 5394 2694
rect 5450 2692 5474 2694
rect 5530 2692 5536 2694
rect 5228 2683 5536 2692
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5172 2576 5224 2582
rect 5172 2518 5224 2524
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 3036 2204 3344 2213
rect 3036 2202 3042 2204
rect 3098 2202 3122 2204
rect 3178 2202 3202 2204
rect 3258 2202 3282 2204
rect 3338 2202 3344 2204
rect 3098 2150 3100 2202
rect 3280 2150 3282 2202
rect 3036 2148 3042 2150
rect 3098 2148 3122 2150
rect 3178 2148 3202 2150
rect 3258 2148 3282 2150
rect 3338 2148 3344 2150
rect 3036 2139 3344 2148
rect 4540 800 4568 2246
rect 5184 800 5212 2518
rect 5736 2514 5764 2746
rect 7024 2514 7052 2994
rect 7944 2650 7972 2994
rect 8080 2748 8388 2757
rect 8080 2746 8086 2748
rect 8142 2746 8166 2748
rect 8222 2746 8246 2748
rect 8302 2746 8326 2748
rect 8382 2746 8388 2748
rect 8142 2694 8144 2746
rect 8324 2694 8326 2746
rect 8080 2692 8086 2694
rect 8142 2692 8166 2694
rect 8222 2692 8246 2694
rect 8302 2692 8326 2694
rect 8382 2692 8388 2694
rect 8080 2683 8388 2692
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 8496 2446 8524 3878
rect 8740 3292 9048 3301
rect 8740 3290 8746 3292
rect 8802 3290 8826 3292
rect 8882 3290 8906 3292
rect 8962 3290 8986 3292
rect 9042 3290 9048 3292
rect 8802 3238 8804 3290
rect 8984 3238 8986 3290
rect 8740 3236 8746 3238
rect 8802 3236 8826 3238
rect 8882 3236 8906 3238
rect 8962 3236 8986 3238
rect 9042 3236 9048 3238
rect 8740 3227 9048 3236
rect 9232 2854 9260 3878
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 9324 3466 9352 3606
rect 9416 3534 9444 4558
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9324 3194 9352 3402
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9416 2514 9444 3470
rect 9784 3058 9812 3538
rect 9876 3126 9904 6151
rect 10152 5642 10180 7346
rect 10244 6322 10272 9030
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10336 8498 10364 8842
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10336 8362 10364 8434
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10520 8294 10548 8842
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10428 7546 10456 7822
rect 10520 7818 10548 8230
rect 10508 7812 10560 7818
rect 10508 7754 10560 7760
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10520 7478 10548 7754
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10244 5710 10272 6258
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5846 10456 6190
rect 10520 5914 10548 6802
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10416 5840 10468 5846
rect 10416 5782 10468 5788
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10140 5636 10192 5642
rect 10140 5578 10192 5584
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9968 4622 9996 5170
rect 10152 4826 10180 5170
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 9956 4616 10008 4622
rect 9956 4558 10008 4564
rect 9968 3670 9996 4558
rect 10244 4486 10272 5646
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10244 4282 10272 4422
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 9968 3074 9996 3606
rect 10060 3534 10088 3946
rect 10152 3534 10180 4150
rect 10336 4146 10364 4694
rect 10428 4690 10456 5782
rect 10508 5704 10560 5710
rect 10612 5692 10640 10798
rect 10692 10668 10744 10674
rect 10692 10610 10744 10616
rect 10704 10062 10732 10610
rect 10796 10606 10824 11086
rect 10876 11076 10928 11082
rect 10876 11018 10928 11024
rect 10888 10742 10916 11018
rect 11592 10908 11900 10917
rect 11592 10906 11598 10908
rect 11654 10906 11678 10908
rect 11734 10906 11758 10908
rect 11814 10906 11838 10908
rect 11894 10906 11900 10908
rect 11654 10854 11656 10906
rect 11836 10854 11838 10906
rect 11592 10852 11598 10854
rect 11654 10852 11678 10854
rect 11734 10852 11758 10854
rect 11814 10852 11838 10854
rect 11894 10852 11900 10854
rect 11592 10843 11900 10852
rect 10876 10736 10928 10742
rect 10876 10678 10928 10684
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 10796 10062 10824 10406
rect 10932 10364 11240 10373
rect 10932 10362 10938 10364
rect 10994 10362 11018 10364
rect 11074 10362 11098 10364
rect 11154 10362 11178 10364
rect 11234 10362 11240 10364
rect 10994 10310 10996 10362
rect 11176 10310 11178 10362
rect 10932 10308 10938 10310
rect 10994 10308 11018 10310
rect 11074 10308 11098 10310
rect 11154 10308 11178 10310
rect 11234 10308 11240 10310
rect 10932 10299 11240 10308
rect 11428 10124 11480 10130
rect 11428 10066 11480 10072
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10784 10056 10836 10062
rect 10784 9998 10836 10004
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 10932 9276 11240 9285
rect 10932 9274 10938 9276
rect 10994 9274 11018 9276
rect 11074 9274 11098 9276
rect 11154 9274 11178 9276
rect 11234 9274 11240 9276
rect 10994 9222 10996 9274
rect 11176 9222 11178 9274
rect 10932 9220 10938 9222
rect 10994 9220 11018 9222
rect 11074 9220 11098 9222
rect 11154 9220 11178 9222
rect 11234 9220 11240 9222
rect 10932 9211 11240 9220
rect 11348 9058 11376 9862
rect 10692 9036 10744 9042
rect 10692 8978 10744 8984
rect 11256 9030 11376 9058
rect 10704 8498 10732 8978
rect 11256 8906 11284 9030
rect 11336 8968 11388 8974
rect 11336 8910 11388 8916
rect 11244 8900 11296 8906
rect 11244 8842 11296 8848
rect 11348 8634 11376 8910
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10796 8090 10824 8366
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 10932 8188 11240 8197
rect 10932 8186 10938 8188
rect 10994 8186 11018 8188
rect 11074 8186 11098 8188
rect 11154 8186 11178 8188
rect 11234 8186 11240 8188
rect 10994 8134 10996 8186
rect 11176 8134 11178 8186
rect 10932 8132 10938 8134
rect 10994 8132 11018 8134
rect 11074 8132 11098 8134
rect 11154 8132 11178 8134
rect 11234 8132 11240 8134
rect 10932 8123 11240 8132
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 10980 7410 11008 7958
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10704 6798 10732 7346
rect 11348 7342 11376 8298
rect 11440 7834 11468 10066
rect 11592 9820 11900 9829
rect 11592 9818 11598 9820
rect 11654 9818 11678 9820
rect 11734 9818 11758 9820
rect 11814 9818 11838 9820
rect 11894 9818 11900 9820
rect 11654 9766 11656 9818
rect 11836 9766 11838 9818
rect 11592 9764 11598 9766
rect 11654 9764 11678 9766
rect 11734 9764 11758 9766
rect 11814 9764 11838 9766
rect 11894 9764 11900 9766
rect 11592 9755 11900 9764
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11532 8634 11560 8774
rect 11592 8732 11900 8741
rect 11592 8730 11598 8732
rect 11654 8730 11678 8732
rect 11734 8730 11758 8732
rect 11814 8730 11838 8732
rect 11894 8730 11900 8732
rect 11654 8678 11656 8730
rect 11836 8678 11838 8730
rect 11592 8676 11598 8678
rect 11654 8676 11678 8678
rect 11734 8676 11758 8678
rect 11814 8676 11838 8678
rect 11894 8676 11900 8678
rect 11592 8667 11900 8676
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11808 7886 11836 8434
rect 11796 7880 11848 7886
rect 11440 7806 11560 7834
rect 11796 7822 11848 7828
rect 11428 7744 11480 7750
rect 11428 7686 11480 7692
rect 11440 7410 11468 7686
rect 11532 7546 11560 7806
rect 11592 7644 11900 7653
rect 11592 7642 11598 7644
rect 11654 7642 11678 7644
rect 11734 7642 11758 7644
rect 11814 7642 11838 7644
rect 11894 7642 11900 7644
rect 11654 7590 11656 7642
rect 11836 7590 11838 7642
rect 11592 7588 11598 7590
rect 11654 7588 11678 7590
rect 11734 7588 11758 7590
rect 11814 7588 11838 7590
rect 11894 7588 11900 7590
rect 11592 7579 11900 7588
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11992 7410 12020 10406
rect 12070 8936 12126 8945
rect 12070 8871 12126 8880
rect 12084 8838 12112 8871
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11336 7336 11388 7342
rect 10796 7274 10916 7290
rect 11336 7278 11388 7284
rect 10796 7268 10928 7274
rect 10796 7262 10876 7268
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10796 6390 10824 7262
rect 10876 7210 10928 7216
rect 10932 7100 11240 7109
rect 10932 7098 10938 7100
rect 10994 7098 11018 7100
rect 11074 7098 11098 7100
rect 11154 7098 11178 7100
rect 11234 7098 11240 7100
rect 10994 7046 10996 7098
rect 11176 7046 11178 7098
rect 10932 7044 10938 7046
rect 10994 7044 11018 7046
rect 11074 7044 11098 7046
rect 11154 7044 11178 7046
rect 11234 7044 11240 7046
rect 10932 7035 11240 7044
rect 11348 6798 11376 7278
rect 11440 6866 11468 7346
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10980 6458 11008 6598
rect 11532 6458 11560 7346
rect 11980 6928 12032 6934
rect 11980 6870 12032 6876
rect 12162 6896 12218 6905
rect 11592 6556 11900 6565
rect 11592 6554 11598 6556
rect 11654 6554 11678 6556
rect 11734 6554 11758 6556
rect 11814 6554 11838 6556
rect 11894 6554 11900 6556
rect 11654 6502 11656 6554
rect 11836 6502 11838 6554
rect 11592 6500 11598 6502
rect 11654 6500 11678 6502
rect 11734 6500 11758 6502
rect 11814 6500 11838 6502
rect 11894 6500 11900 6502
rect 11592 6491 11900 6500
rect 10968 6452 11020 6458
rect 10968 6394 11020 6400
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 11992 6390 12020 6870
rect 12162 6831 12164 6840
rect 12216 6831 12218 6840
rect 12164 6802 12216 6808
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11610 6216 11666 6225
rect 11336 6180 11388 6186
rect 11610 6151 11612 6160
rect 11336 6122 11388 6128
rect 11664 6151 11666 6160
rect 11612 6122 11664 6128
rect 10932 6012 11240 6021
rect 10932 6010 10938 6012
rect 10994 6010 11018 6012
rect 11074 6010 11098 6012
rect 11154 6010 11178 6012
rect 11234 6010 11240 6012
rect 10994 5958 10996 6010
rect 11176 5958 11178 6010
rect 10932 5956 10938 5958
rect 10994 5956 11018 5958
rect 11074 5956 11098 5958
rect 11154 5956 11178 5958
rect 11234 5956 11240 5958
rect 10932 5947 11240 5956
rect 11348 5778 11376 6122
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 10784 5704 10836 5710
rect 10612 5664 10784 5692
rect 10508 5646 10560 5652
rect 10784 5646 10836 5652
rect 10520 5370 10548 5646
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10704 4826 10732 5510
rect 11440 5302 11468 6054
rect 11592 5468 11900 5477
rect 11592 5466 11598 5468
rect 11654 5466 11678 5468
rect 11734 5466 11758 5468
rect 11814 5466 11838 5468
rect 11894 5466 11900 5468
rect 11654 5414 11656 5466
rect 11836 5414 11838 5466
rect 11592 5412 11598 5414
rect 11654 5412 11678 5414
rect 11734 5412 11758 5414
rect 11814 5412 11838 5414
rect 11894 5412 11900 5414
rect 11592 5403 11900 5412
rect 11428 5296 11480 5302
rect 11428 5238 11480 5244
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 10932 4924 11240 4933
rect 10932 4922 10938 4924
rect 10994 4922 11018 4924
rect 11074 4922 11098 4924
rect 11154 4922 11178 4924
rect 11234 4922 11240 4924
rect 10994 4870 10996 4922
rect 11176 4870 11178 4922
rect 10932 4868 10938 4870
rect 10994 4868 11018 4870
rect 11074 4868 11098 4870
rect 11154 4868 11178 4870
rect 11234 4868 11240 4870
rect 10932 4859 11240 4868
rect 11716 4865 11744 4966
rect 11702 4856 11758 4865
rect 10692 4820 10744 4826
rect 11992 4826 12020 6326
rect 12070 6216 12126 6225
rect 12070 6151 12126 6160
rect 12084 5370 12112 6151
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12176 5545 12204 5646
rect 12162 5536 12218 5545
rect 12162 5471 12218 5480
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11702 4791 11758 4800
rect 11980 4820 12032 4826
rect 10692 4762 10744 4768
rect 11980 4762 12032 4768
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 10428 4214 10456 4626
rect 10416 4208 10468 4214
rect 10416 4150 10468 4156
rect 10692 4208 10744 4214
rect 10692 4150 10744 4156
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10336 3942 10364 4082
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3534 10364 3878
rect 10428 3738 10456 3946
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 10060 3194 10088 3470
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 9772 3052 9824 3058
rect 9968 3046 10088 3074
rect 9772 2994 9824 3000
rect 10060 2854 10088 3046
rect 10152 2990 10180 3470
rect 10428 3058 10456 3674
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10612 2990 10640 4082
rect 10704 3466 10732 4150
rect 10980 4026 11008 4626
rect 11520 4548 11572 4554
rect 11520 4490 11572 4496
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 11164 4214 11192 4422
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11532 4078 11560 4490
rect 11592 4380 11900 4389
rect 11592 4378 11598 4380
rect 11654 4378 11678 4380
rect 11734 4378 11758 4380
rect 11814 4378 11838 4380
rect 11894 4378 11900 4380
rect 11654 4326 11656 4378
rect 11836 4326 11838 4378
rect 11592 4324 11598 4326
rect 11654 4324 11678 4326
rect 11734 4324 11758 4326
rect 11814 4324 11838 4326
rect 11894 4324 11900 4326
rect 11592 4315 11900 4324
rect 10796 4010 11008 4026
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 10784 4004 11008 4010
rect 10836 3998 11008 4004
rect 10784 3946 10836 3952
rect 10692 3460 10744 3466
rect 10692 3402 10744 3408
rect 10796 3194 10824 3946
rect 10932 3836 11240 3845
rect 10932 3834 10938 3836
rect 10994 3834 11018 3836
rect 11074 3834 11098 3836
rect 11154 3834 11178 3836
rect 11234 3834 11240 3836
rect 10994 3782 10996 3834
rect 11176 3782 11178 3834
rect 10932 3780 10938 3782
rect 10994 3780 11018 3782
rect 11074 3780 11098 3782
rect 11154 3780 11178 3782
rect 11234 3780 11240 3782
rect 10932 3771 11240 3780
rect 11592 3292 11900 3301
rect 11592 3290 11598 3292
rect 11654 3290 11678 3292
rect 11734 3290 11758 3292
rect 11814 3290 11838 3292
rect 11894 3290 11900 3292
rect 11654 3238 11656 3290
rect 11836 3238 11838 3290
rect 11592 3236 11598 3238
rect 11654 3236 11678 3238
rect 11734 3236 11758 3238
rect 11814 3236 11838 3238
rect 11894 3236 11900 3238
rect 11592 3227 11900 3236
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2650 10088 2790
rect 10932 2748 11240 2757
rect 10932 2746 10938 2748
rect 10994 2746 11018 2748
rect 11074 2746 11098 2748
rect 11154 2746 11178 2748
rect 11234 2746 11240 2748
rect 10994 2694 10996 2746
rect 11176 2694 11178 2746
rect 10932 2692 10938 2694
rect 10994 2692 11018 2694
rect 11074 2692 11098 2694
rect 11154 2692 11178 2694
rect 11234 2692 11240 2694
rect 10932 2683 11240 2692
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 5828 800 5856 2382
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 5888 2204 6196 2213
rect 5888 2202 5894 2204
rect 5950 2202 5974 2204
rect 6030 2202 6054 2204
rect 6110 2202 6134 2204
rect 6190 2202 6196 2204
rect 5950 2150 5952 2202
rect 6132 2150 6134 2202
rect 5888 2148 5894 2150
rect 5950 2148 5974 2150
rect 6030 2148 6054 2150
rect 6110 2148 6134 2150
rect 6190 2148 6196 2150
rect 5888 2139 6196 2148
rect 6472 800 6500 2314
rect 7116 800 7144 2382
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 7760 800 7788 2246
rect 8404 800 8432 2246
rect 8740 2204 9048 2213
rect 8740 2202 8746 2204
rect 8802 2202 8826 2204
rect 8882 2202 8906 2204
rect 8962 2202 8986 2204
rect 9042 2202 9048 2204
rect 8802 2150 8804 2202
rect 8984 2150 8986 2202
rect 8740 2148 8746 2150
rect 8802 2148 8826 2150
rect 8882 2148 8906 2150
rect 8962 2148 8986 2150
rect 9042 2148 9048 2150
rect 8740 2139 9048 2148
rect 9140 1306 9168 2382
rect 9048 1278 9168 1306
rect 9048 800 9076 1278
rect 9692 800 9720 2382
rect 11592 2204 11900 2213
rect 11592 2202 11598 2204
rect 11654 2202 11678 2204
rect 11734 2202 11758 2204
rect 11814 2202 11838 2204
rect 11894 2202 11900 2204
rect 11654 2150 11656 2202
rect 11836 2150 11838 2202
rect 11592 2148 11598 2150
rect 11654 2148 11678 2150
rect 11734 2148 11758 2150
rect 11814 2148 11838 2150
rect 11894 2148 11900 2150
rect 11592 2139 11900 2148
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
<< via2 >>
rect 2382 13626 2438 13628
rect 2462 13626 2518 13628
rect 2542 13626 2598 13628
rect 2622 13626 2678 13628
rect 2382 13574 2428 13626
rect 2428 13574 2438 13626
rect 2462 13574 2492 13626
rect 2492 13574 2504 13626
rect 2504 13574 2518 13626
rect 2542 13574 2556 13626
rect 2556 13574 2568 13626
rect 2568 13574 2598 13626
rect 2622 13574 2632 13626
rect 2632 13574 2678 13626
rect 2382 13572 2438 13574
rect 2462 13572 2518 13574
rect 2542 13572 2598 13574
rect 2622 13572 2678 13574
rect 5234 13626 5290 13628
rect 5314 13626 5370 13628
rect 5394 13626 5450 13628
rect 5474 13626 5530 13628
rect 5234 13574 5280 13626
rect 5280 13574 5290 13626
rect 5314 13574 5344 13626
rect 5344 13574 5356 13626
rect 5356 13574 5370 13626
rect 5394 13574 5408 13626
rect 5408 13574 5420 13626
rect 5420 13574 5450 13626
rect 5474 13574 5484 13626
rect 5484 13574 5530 13626
rect 5234 13572 5290 13574
rect 5314 13572 5370 13574
rect 5394 13572 5450 13574
rect 5474 13572 5530 13574
rect 8086 13626 8142 13628
rect 8166 13626 8222 13628
rect 8246 13626 8302 13628
rect 8326 13626 8382 13628
rect 8086 13574 8132 13626
rect 8132 13574 8142 13626
rect 8166 13574 8196 13626
rect 8196 13574 8208 13626
rect 8208 13574 8222 13626
rect 8246 13574 8260 13626
rect 8260 13574 8272 13626
rect 8272 13574 8302 13626
rect 8326 13574 8336 13626
rect 8336 13574 8382 13626
rect 8086 13572 8142 13574
rect 8166 13572 8222 13574
rect 8246 13572 8302 13574
rect 8326 13572 8382 13574
rect 10938 13626 10994 13628
rect 11018 13626 11074 13628
rect 11098 13626 11154 13628
rect 11178 13626 11234 13628
rect 10938 13574 10984 13626
rect 10984 13574 10994 13626
rect 11018 13574 11048 13626
rect 11048 13574 11060 13626
rect 11060 13574 11074 13626
rect 11098 13574 11112 13626
rect 11112 13574 11124 13626
rect 11124 13574 11154 13626
rect 11178 13574 11188 13626
rect 11188 13574 11234 13626
rect 10938 13572 10994 13574
rect 11018 13572 11074 13574
rect 11098 13572 11154 13574
rect 11178 13572 11234 13574
rect 3042 13082 3098 13084
rect 3122 13082 3178 13084
rect 3202 13082 3258 13084
rect 3282 13082 3338 13084
rect 3042 13030 3088 13082
rect 3088 13030 3098 13082
rect 3122 13030 3152 13082
rect 3152 13030 3164 13082
rect 3164 13030 3178 13082
rect 3202 13030 3216 13082
rect 3216 13030 3228 13082
rect 3228 13030 3258 13082
rect 3282 13030 3292 13082
rect 3292 13030 3338 13082
rect 3042 13028 3098 13030
rect 3122 13028 3178 13030
rect 3202 13028 3258 13030
rect 3282 13028 3338 13030
rect 1398 12280 1454 12336
rect 1030 11600 1086 11656
rect 2382 12538 2438 12540
rect 2462 12538 2518 12540
rect 2542 12538 2598 12540
rect 2622 12538 2678 12540
rect 2382 12486 2428 12538
rect 2428 12486 2438 12538
rect 2462 12486 2492 12538
rect 2492 12486 2504 12538
rect 2504 12486 2518 12538
rect 2542 12486 2556 12538
rect 2556 12486 2568 12538
rect 2568 12486 2598 12538
rect 2622 12486 2632 12538
rect 2632 12486 2678 12538
rect 2382 12484 2438 12486
rect 2462 12484 2518 12486
rect 2542 12484 2598 12486
rect 2622 12484 2678 12486
rect 3042 11994 3098 11996
rect 3122 11994 3178 11996
rect 3202 11994 3258 11996
rect 3282 11994 3338 11996
rect 3042 11942 3088 11994
rect 3088 11942 3098 11994
rect 3122 11942 3152 11994
rect 3152 11942 3164 11994
rect 3164 11942 3178 11994
rect 3202 11942 3216 11994
rect 3216 11942 3228 11994
rect 3228 11942 3258 11994
rect 3282 11942 3292 11994
rect 3292 11942 3338 11994
rect 3042 11940 3098 11942
rect 3122 11940 3178 11942
rect 3202 11940 3258 11942
rect 3282 11940 3338 11942
rect 2382 11450 2438 11452
rect 2462 11450 2518 11452
rect 2542 11450 2598 11452
rect 2622 11450 2678 11452
rect 2382 11398 2428 11450
rect 2428 11398 2438 11450
rect 2462 11398 2492 11450
rect 2492 11398 2504 11450
rect 2504 11398 2518 11450
rect 2542 11398 2556 11450
rect 2556 11398 2568 11450
rect 2568 11398 2598 11450
rect 2622 11398 2632 11450
rect 2632 11398 2678 11450
rect 2382 11396 2438 11398
rect 2462 11396 2518 11398
rect 2542 11396 2598 11398
rect 2622 11396 2678 11398
rect 1398 10920 1454 10976
rect 3042 10906 3098 10908
rect 3122 10906 3178 10908
rect 3202 10906 3258 10908
rect 3282 10906 3338 10908
rect 3042 10854 3088 10906
rect 3088 10854 3098 10906
rect 3122 10854 3152 10906
rect 3152 10854 3164 10906
rect 3164 10854 3178 10906
rect 3202 10854 3216 10906
rect 3216 10854 3228 10906
rect 3228 10854 3258 10906
rect 3282 10854 3292 10906
rect 3292 10854 3338 10906
rect 3042 10852 3098 10854
rect 3122 10852 3178 10854
rect 3202 10852 3258 10854
rect 3282 10852 3338 10854
rect 1674 9560 1730 9616
rect 1490 9036 1546 9072
rect 1490 9016 1492 9036
rect 1492 9016 1544 9036
rect 1544 9016 1546 9036
rect 1490 8880 1546 8936
rect 1306 8200 1362 8256
rect 938 7520 994 7576
rect 2382 10362 2438 10364
rect 2462 10362 2518 10364
rect 2542 10362 2598 10364
rect 2622 10362 2678 10364
rect 2382 10310 2428 10362
rect 2428 10310 2438 10362
rect 2462 10310 2492 10362
rect 2492 10310 2504 10362
rect 2504 10310 2518 10362
rect 2542 10310 2556 10362
rect 2556 10310 2568 10362
rect 2568 10310 2598 10362
rect 2622 10310 2632 10362
rect 2632 10310 2678 10362
rect 2382 10308 2438 10310
rect 2462 10308 2518 10310
rect 2542 10308 2598 10310
rect 2622 10308 2678 10310
rect 4526 12180 4528 12200
rect 4528 12180 4580 12200
rect 4580 12180 4582 12200
rect 4526 12144 4582 12180
rect 3042 9818 3098 9820
rect 3122 9818 3178 9820
rect 3202 9818 3258 9820
rect 3282 9818 3338 9820
rect 3042 9766 3088 9818
rect 3088 9766 3098 9818
rect 3122 9766 3152 9818
rect 3152 9766 3164 9818
rect 3164 9766 3178 9818
rect 3202 9766 3216 9818
rect 3216 9766 3228 9818
rect 3228 9766 3258 9818
rect 3282 9766 3292 9818
rect 3292 9766 3338 9818
rect 3042 9764 3098 9766
rect 3122 9764 3178 9766
rect 3202 9764 3258 9766
rect 3282 9764 3338 9766
rect 2594 9460 2596 9480
rect 2596 9460 2648 9480
rect 2648 9460 2650 9480
rect 2594 9424 2650 9460
rect 2382 9274 2438 9276
rect 2462 9274 2518 9276
rect 2542 9274 2598 9276
rect 2622 9274 2678 9276
rect 2382 9222 2428 9274
rect 2428 9222 2438 9274
rect 2462 9222 2492 9274
rect 2492 9222 2504 9274
rect 2504 9222 2518 9274
rect 2542 9222 2556 9274
rect 2556 9222 2568 9274
rect 2568 9222 2598 9274
rect 2622 9222 2632 9274
rect 2632 9222 2678 9274
rect 2382 9220 2438 9222
rect 2462 9220 2518 9222
rect 2542 9220 2598 9222
rect 2622 9220 2678 9222
rect 2226 9016 2282 9072
rect 2594 8472 2650 8528
rect 3146 9580 3202 9616
rect 3146 9560 3148 9580
rect 3148 9560 3200 9580
rect 3200 9560 3202 9580
rect 3042 8730 3098 8732
rect 3122 8730 3178 8732
rect 3202 8730 3258 8732
rect 3282 8730 3338 8732
rect 3042 8678 3088 8730
rect 3088 8678 3098 8730
rect 3122 8678 3152 8730
rect 3152 8678 3164 8730
rect 3164 8678 3178 8730
rect 3202 8678 3216 8730
rect 3216 8678 3228 8730
rect 3228 8678 3258 8730
rect 3282 8678 3292 8730
rect 3292 8678 3338 8730
rect 3042 8676 3098 8678
rect 3122 8676 3178 8678
rect 3202 8676 3258 8678
rect 3282 8676 3338 8678
rect 3146 8336 3202 8392
rect 2382 8186 2438 8188
rect 2462 8186 2518 8188
rect 2542 8186 2598 8188
rect 2622 8186 2678 8188
rect 2382 8134 2428 8186
rect 2428 8134 2438 8186
rect 2462 8134 2492 8186
rect 2492 8134 2504 8186
rect 2504 8134 2518 8186
rect 2542 8134 2556 8186
rect 2556 8134 2568 8186
rect 2568 8134 2598 8186
rect 2622 8134 2632 8186
rect 2632 8134 2678 8186
rect 2382 8132 2438 8134
rect 2462 8132 2518 8134
rect 2542 8132 2598 8134
rect 2622 8132 2678 8134
rect 1490 6840 1546 6896
rect 846 6024 902 6080
rect 1490 5480 1546 5536
rect 3042 7642 3098 7644
rect 3122 7642 3178 7644
rect 3202 7642 3258 7644
rect 3282 7642 3338 7644
rect 3042 7590 3088 7642
rect 3088 7590 3098 7642
rect 3122 7590 3152 7642
rect 3152 7590 3164 7642
rect 3164 7590 3178 7642
rect 3202 7590 3216 7642
rect 3216 7590 3228 7642
rect 3228 7590 3258 7642
rect 3282 7590 3292 7642
rect 3292 7590 3338 7642
rect 3042 7588 3098 7590
rect 3122 7588 3178 7590
rect 3202 7588 3258 7590
rect 3282 7588 3338 7590
rect 2382 7098 2438 7100
rect 2462 7098 2518 7100
rect 2542 7098 2598 7100
rect 2622 7098 2678 7100
rect 2382 7046 2428 7098
rect 2428 7046 2438 7098
rect 2462 7046 2492 7098
rect 2492 7046 2504 7098
rect 2504 7046 2518 7098
rect 2542 7046 2556 7098
rect 2556 7046 2568 7098
rect 2568 7046 2598 7098
rect 2622 7046 2632 7098
rect 2632 7046 2678 7098
rect 2382 7044 2438 7046
rect 2462 7044 2518 7046
rect 2542 7044 2598 7046
rect 2622 7044 2678 7046
rect 3042 6554 3098 6556
rect 3122 6554 3178 6556
rect 3202 6554 3258 6556
rect 3282 6554 3338 6556
rect 3042 6502 3088 6554
rect 3088 6502 3098 6554
rect 3122 6502 3152 6554
rect 3152 6502 3164 6554
rect 3164 6502 3178 6554
rect 3202 6502 3216 6554
rect 3216 6502 3228 6554
rect 3228 6502 3258 6554
rect 3282 6502 3292 6554
rect 3292 6502 3338 6554
rect 3042 6500 3098 6502
rect 3122 6500 3178 6502
rect 3202 6500 3258 6502
rect 3282 6500 3338 6502
rect 2382 6010 2438 6012
rect 2462 6010 2518 6012
rect 2542 6010 2598 6012
rect 2622 6010 2678 6012
rect 2382 5958 2428 6010
rect 2428 5958 2438 6010
rect 2462 5958 2492 6010
rect 2492 5958 2504 6010
rect 2504 5958 2518 6010
rect 2542 5958 2556 6010
rect 2556 5958 2568 6010
rect 2568 5958 2598 6010
rect 2622 5958 2632 6010
rect 2632 5958 2678 6010
rect 2382 5956 2438 5958
rect 2462 5956 2518 5958
rect 2542 5956 2598 5958
rect 2622 5956 2678 5958
rect 5894 13082 5950 13084
rect 5974 13082 6030 13084
rect 6054 13082 6110 13084
rect 6134 13082 6190 13084
rect 5894 13030 5940 13082
rect 5940 13030 5950 13082
rect 5974 13030 6004 13082
rect 6004 13030 6016 13082
rect 6016 13030 6030 13082
rect 6054 13030 6068 13082
rect 6068 13030 6080 13082
rect 6080 13030 6110 13082
rect 6134 13030 6144 13082
rect 6144 13030 6190 13082
rect 5894 13028 5950 13030
rect 5974 13028 6030 13030
rect 6054 13028 6110 13030
rect 6134 13028 6190 13030
rect 5234 12538 5290 12540
rect 5314 12538 5370 12540
rect 5394 12538 5450 12540
rect 5474 12538 5530 12540
rect 5234 12486 5280 12538
rect 5280 12486 5290 12538
rect 5314 12486 5344 12538
rect 5344 12486 5356 12538
rect 5356 12486 5370 12538
rect 5394 12486 5408 12538
rect 5408 12486 5420 12538
rect 5420 12486 5450 12538
rect 5474 12486 5484 12538
rect 5484 12486 5530 12538
rect 5234 12484 5290 12486
rect 5314 12484 5370 12486
rect 5394 12484 5450 12486
rect 5474 12484 5530 12486
rect 4250 9016 4306 9072
rect 5262 12144 5318 12200
rect 5894 11994 5950 11996
rect 5974 11994 6030 11996
rect 6054 11994 6110 11996
rect 6134 11994 6190 11996
rect 5894 11942 5940 11994
rect 5940 11942 5950 11994
rect 5974 11942 6004 11994
rect 6004 11942 6016 11994
rect 6016 11942 6030 11994
rect 6054 11942 6068 11994
rect 6068 11942 6080 11994
rect 6080 11942 6110 11994
rect 6134 11942 6144 11994
rect 6144 11942 6190 11994
rect 5894 11940 5950 11942
rect 5974 11940 6030 11942
rect 6054 11940 6110 11942
rect 6134 11940 6190 11942
rect 5234 11450 5290 11452
rect 5314 11450 5370 11452
rect 5394 11450 5450 11452
rect 5474 11450 5530 11452
rect 5234 11398 5280 11450
rect 5280 11398 5290 11450
rect 5314 11398 5344 11450
rect 5344 11398 5356 11450
rect 5356 11398 5370 11450
rect 5394 11398 5408 11450
rect 5408 11398 5420 11450
rect 5420 11398 5450 11450
rect 5474 11398 5484 11450
rect 5484 11398 5530 11450
rect 5234 11396 5290 11398
rect 5314 11396 5370 11398
rect 5394 11396 5450 11398
rect 5474 11396 5530 11398
rect 8746 13082 8802 13084
rect 8826 13082 8882 13084
rect 8906 13082 8962 13084
rect 8986 13082 9042 13084
rect 8746 13030 8792 13082
rect 8792 13030 8802 13082
rect 8826 13030 8856 13082
rect 8856 13030 8868 13082
rect 8868 13030 8882 13082
rect 8906 13030 8920 13082
rect 8920 13030 8932 13082
rect 8932 13030 8962 13082
rect 8986 13030 8996 13082
rect 8996 13030 9042 13082
rect 8746 13028 8802 13030
rect 8826 13028 8882 13030
rect 8906 13028 8962 13030
rect 8986 13028 9042 13030
rect 11598 13082 11654 13084
rect 11678 13082 11734 13084
rect 11758 13082 11814 13084
rect 11838 13082 11894 13084
rect 11598 13030 11644 13082
rect 11644 13030 11654 13082
rect 11678 13030 11708 13082
rect 11708 13030 11720 13082
rect 11720 13030 11734 13082
rect 11758 13030 11772 13082
rect 11772 13030 11784 13082
rect 11784 13030 11814 13082
rect 11838 13030 11848 13082
rect 11848 13030 11894 13082
rect 11598 13028 11654 13030
rect 11678 13028 11734 13030
rect 11758 13028 11814 13030
rect 11838 13028 11894 13030
rect 8086 12538 8142 12540
rect 8166 12538 8222 12540
rect 8246 12538 8302 12540
rect 8326 12538 8382 12540
rect 8086 12486 8132 12538
rect 8132 12486 8142 12538
rect 8166 12486 8196 12538
rect 8196 12486 8208 12538
rect 8208 12486 8222 12538
rect 8246 12486 8260 12538
rect 8260 12486 8272 12538
rect 8272 12486 8302 12538
rect 8326 12486 8336 12538
rect 8336 12486 8382 12538
rect 8086 12484 8142 12486
rect 8166 12484 8222 12486
rect 8246 12484 8302 12486
rect 8326 12484 8382 12486
rect 8746 11994 8802 11996
rect 8826 11994 8882 11996
rect 8906 11994 8962 11996
rect 8986 11994 9042 11996
rect 8746 11942 8792 11994
rect 8792 11942 8802 11994
rect 8826 11942 8856 11994
rect 8856 11942 8868 11994
rect 8868 11942 8882 11994
rect 8906 11942 8920 11994
rect 8920 11942 8932 11994
rect 8932 11942 8962 11994
rect 8986 11942 8996 11994
rect 8996 11942 9042 11994
rect 8746 11940 8802 11942
rect 8826 11940 8882 11942
rect 8906 11940 8962 11942
rect 8986 11940 9042 11942
rect 5894 10906 5950 10908
rect 5974 10906 6030 10908
rect 6054 10906 6110 10908
rect 6134 10906 6190 10908
rect 5894 10854 5940 10906
rect 5940 10854 5950 10906
rect 5974 10854 6004 10906
rect 6004 10854 6016 10906
rect 6016 10854 6030 10906
rect 6054 10854 6068 10906
rect 6068 10854 6080 10906
rect 6080 10854 6110 10906
rect 6134 10854 6144 10906
rect 6144 10854 6190 10906
rect 5894 10852 5950 10854
rect 5974 10852 6030 10854
rect 6054 10852 6110 10854
rect 6134 10852 6190 10854
rect 4526 8356 4582 8392
rect 4526 8336 4528 8356
rect 4528 8336 4580 8356
rect 4580 8336 4582 8356
rect 846 4936 902 4992
rect 2382 4922 2438 4924
rect 2462 4922 2518 4924
rect 2542 4922 2598 4924
rect 2622 4922 2678 4924
rect 2382 4870 2428 4922
rect 2428 4870 2438 4922
rect 2462 4870 2492 4922
rect 2492 4870 2504 4922
rect 2504 4870 2518 4922
rect 2542 4870 2556 4922
rect 2556 4870 2568 4922
rect 2568 4870 2598 4922
rect 2622 4870 2632 4922
rect 2632 4870 2678 4922
rect 2382 4868 2438 4870
rect 2462 4868 2518 4870
rect 2542 4868 2598 4870
rect 2622 4868 2678 4870
rect 3042 5466 3098 5468
rect 3122 5466 3178 5468
rect 3202 5466 3258 5468
rect 3282 5466 3338 5468
rect 3042 5414 3088 5466
rect 3088 5414 3098 5466
rect 3122 5414 3152 5466
rect 3152 5414 3164 5466
rect 3164 5414 3178 5466
rect 3202 5414 3216 5466
rect 3216 5414 3228 5466
rect 3228 5414 3258 5466
rect 3282 5414 3292 5466
rect 3292 5414 3338 5466
rect 3042 5412 3098 5414
rect 3122 5412 3178 5414
rect 3202 5412 3258 5414
rect 3282 5412 3338 5414
rect 4894 8492 4950 8528
rect 4894 8472 4896 8492
rect 4896 8472 4948 8492
rect 4948 8472 4950 8492
rect 5234 10362 5290 10364
rect 5314 10362 5370 10364
rect 5394 10362 5450 10364
rect 5474 10362 5530 10364
rect 5234 10310 5280 10362
rect 5280 10310 5290 10362
rect 5314 10310 5344 10362
rect 5344 10310 5356 10362
rect 5356 10310 5370 10362
rect 5394 10310 5408 10362
rect 5408 10310 5420 10362
rect 5420 10310 5450 10362
rect 5474 10310 5484 10362
rect 5484 10310 5530 10362
rect 5234 10308 5290 10310
rect 5314 10308 5370 10310
rect 5394 10308 5450 10310
rect 5474 10308 5530 10310
rect 8086 11450 8142 11452
rect 8166 11450 8222 11452
rect 8246 11450 8302 11452
rect 8326 11450 8382 11452
rect 8086 11398 8132 11450
rect 8132 11398 8142 11450
rect 8166 11398 8196 11450
rect 8196 11398 8208 11450
rect 8208 11398 8222 11450
rect 8246 11398 8260 11450
rect 8260 11398 8272 11450
rect 8272 11398 8302 11450
rect 8326 11398 8336 11450
rect 8336 11398 8382 11450
rect 8086 11396 8142 11398
rect 8166 11396 8222 11398
rect 8246 11396 8302 11398
rect 8326 11396 8382 11398
rect 7654 11092 7656 11112
rect 7656 11092 7708 11112
rect 7708 11092 7710 11112
rect 7654 11056 7710 11092
rect 8482 11092 8484 11112
rect 8484 11092 8536 11112
rect 8536 11092 8538 11112
rect 5894 9818 5950 9820
rect 5974 9818 6030 9820
rect 6054 9818 6110 9820
rect 6134 9818 6190 9820
rect 5894 9766 5940 9818
rect 5940 9766 5950 9818
rect 5974 9766 6004 9818
rect 6004 9766 6016 9818
rect 6016 9766 6030 9818
rect 6054 9766 6068 9818
rect 6068 9766 6080 9818
rect 6080 9766 6110 9818
rect 6134 9766 6144 9818
rect 6144 9766 6190 9818
rect 5894 9764 5950 9766
rect 5974 9764 6030 9766
rect 6054 9764 6110 9766
rect 6134 9764 6190 9766
rect 5234 9274 5290 9276
rect 5314 9274 5370 9276
rect 5394 9274 5450 9276
rect 5474 9274 5530 9276
rect 5234 9222 5280 9274
rect 5280 9222 5290 9274
rect 5314 9222 5344 9274
rect 5344 9222 5356 9274
rect 5356 9222 5370 9274
rect 5394 9222 5408 9274
rect 5408 9222 5420 9274
rect 5420 9222 5450 9274
rect 5474 9222 5484 9274
rect 5484 9222 5530 9274
rect 5234 9220 5290 9222
rect 5314 9220 5370 9222
rect 5394 9220 5450 9222
rect 5474 9220 5530 9222
rect 5234 8186 5290 8188
rect 5314 8186 5370 8188
rect 5394 8186 5450 8188
rect 5474 8186 5530 8188
rect 5234 8134 5280 8186
rect 5280 8134 5290 8186
rect 5314 8134 5344 8186
rect 5344 8134 5356 8186
rect 5356 8134 5370 8186
rect 5394 8134 5408 8186
rect 5408 8134 5420 8186
rect 5420 8134 5450 8186
rect 5474 8134 5484 8186
rect 5484 8134 5530 8186
rect 5234 8132 5290 8134
rect 5314 8132 5370 8134
rect 5394 8132 5450 8134
rect 5474 8132 5530 8134
rect 4158 5636 4214 5672
rect 4158 5616 4160 5636
rect 4160 5616 4212 5636
rect 4212 5616 4214 5636
rect 3042 4378 3098 4380
rect 3122 4378 3178 4380
rect 3202 4378 3258 4380
rect 3282 4378 3338 4380
rect 3042 4326 3088 4378
rect 3088 4326 3098 4378
rect 3122 4326 3152 4378
rect 3152 4326 3164 4378
rect 3164 4326 3178 4378
rect 3202 4326 3216 4378
rect 3216 4326 3228 4378
rect 3228 4326 3258 4378
rect 3282 4326 3292 4378
rect 3292 4326 3338 4378
rect 3042 4324 3098 4326
rect 3122 4324 3178 4326
rect 3202 4324 3258 4326
rect 3282 4324 3338 4326
rect 2382 3834 2438 3836
rect 2462 3834 2518 3836
rect 2542 3834 2598 3836
rect 2622 3834 2678 3836
rect 2382 3782 2428 3834
rect 2428 3782 2438 3834
rect 2462 3782 2492 3834
rect 2492 3782 2504 3834
rect 2504 3782 2518 3834
rect 2542 3782 2556 3834
rect 2556 3782 2568 3834
rect 2568 3782 2598 3834
rect 2622 3782 2632 3834
rect 2632 3782 2678 3834
rect 2382 3780 2438 3782
rect 2462 3780 2518 3782
rect 2542 3780 2598 3782
rect 2622 3780 2678 3782
rect 3042 3290 3098 3292
rect 3122 3290 3178 3292
rect 3202 3290 3258 3292
rect 3282 3290 3338 3292
rect 3042 3238 3088 3290
rect 3088 3238 3098 3290
rect 3122 3238 3152 3290
rect 3152 3238 3164 3290
rect 3164 3238 3178 3290
rect 3202 3238 3216 3290
rect 3216 3238 3228 3290
rect 3228 3238 3258 3290
rect 3282 3238 3292 3290
rect 3292 3238 3338 3290
rect 3042 3236 3098 3238
rect 3122 3236 3178 3238
rect 3202 3236 3258 3238
rect 3282 3236 3338 3238
rect 2382 2746 2438 2748
rect 2462 2746 2518 2748
rect 2542 2746 2598 2748
rect 2622 2746 2678 2748
rect 2382 2694 2428 2746
rect 2428 2694 2438 2746
rect 2462 2694 2492 2746
rect 2492 2694 2504 2746
rect 2504 2694 2518 2746
rect 2542 2694 2556 2746
rect 2556 2694 2568 2746
rect 2568 2694 2598 2746
rect 2622 2694 2632 2746
rect 2632 2694 2678 2746
rect 2382 2692 2438 2694
rect 2462 2692 2518 2694
rect 2542 2692 2598 2694
rect 2622 2692 2678 2694
rect 5234 7098 5290 7100
rect 5314 7098 5370 7100
rect 5394 7098 5450 7100
rect 5474 7098 5530 7100
rect 5234 7046 5280 7098
rect 5280 7046 5290 7098
rect 5314 7046 5344 7098
rect 5344 7046 5356 7098
rect 5356 7046 5370 7098
rect 5394 7046 5408 7098
rect 5408 7046 5420 7098
rect 5420 7046 5450 7098
rect 5474 7046 5484 7098
rect 5484 7046 5530 7098
rect 5234 7044 5290 7046
rect 5314 7044 5370 7046
rect 5394 7044 5450 7046
rect 5474 7044 5530 7046
rect 5894 8730 5950 8732
rect 5974 8730 6030 8732
rect 6054 8730 6110 8732
rect 6134 8730 6190 8732
rect 5894 8678 5940 8730
rect 5940 8678 5950 8730
rect 5974 8678 6004 8730
rect 6004 8678 6016 8730
rect 6016 8678 6030 8730
rect 6054 8678 6068 8730
rect 6068 8678 6080 8730
rect 6080 8678 6110 8730
rect 6134 8678 6144 8730
rect 6144 8678 6190 8730
rect 5894 8676 5950 8678
rect 5974 8676 6030 8678
rect 6054 8676 6110 8678
rect 6134 8676 6190 8678
rect 5894 7642 5950 7644
rect 5974 7642 6030 7644
rect 6054 7642 6110 7644
rect 6134 7642 6190 7644
rect 5894 7590 5940 7642
rect 5940 7590 5950 7642
rect 5974 7590 6004 7642
rect 6004 7590 6016 7642
rect 6016 7590 6030 7642
rect 6054 7590 6068 7642
rect 6068 7590 6080 7642
rect 6080 7590 6110 7642
rect 6134 7590 6144 7642
rect 6144 7590 6190 7642
rect 5894 7588 5950 7590
rect 5974 7588 6030 7590
rect 6054 7588 6110 7590
rect 6134 7588 6190 7590
rect 5894 6554 5950 6556
rect 5974 6554 6030 6556
rect 6054 6554 6110 6556
rect 6134 6554 6190 6556
rect 5894 6502 5940 6554
rect 5940 6502 5950 6554
rect 5974 6502 6004 6554
rect 6004 6502 6016 6554
rect 6016 6502 6030 6554
rect 6054 6502 6068 6554
rect 6068 6502 6080 6554
rect 6080 6502 6110 6554
rect 6134 6502 6144 6554
rect 6144 6502 6190 6554
rect 5894 6500 5950 6502
rect 5974 6500 6030 6502
rect 6054 6500 6110 6502
rect 6134 6500 6190 6502
rect 5234 6010 5290 6012
rect 5314 6010 5370 6012
rect 5394 6010 5450 6012
rect 5474 6010 5530 6012
rect 5234 5958 5280 6010
rect 5280 5958 5290 6010
rect 5314 5958 5344 6010
rect 5344 5958 5356 6010
rect 5356 5958 5370 6010
rect 5394 5958 5408 6010
rect 5408 5958 5420 6010
rect 5420 5958 5450 6010
rect 5474 5958 5484 6010
rect 5484 5958 5530 6010
rect 5234 5956 5290 5958
rect 5314 5956 5370 5958
rect 5394 5956 5450 5958
rect 5474 5956 5530 5958
rect 5998 5652 6000 5672
rect 6000 5652 6052 5672
rect 6052 5652 6054 5672
rect 5234 4922 5290 4924
rect 5314 4922 5370 4924
rect 5394 4922 5450 4924
rect 5474 4922 5530 4924
rect 5234 4870 5280 4922
rect 5280 4870 5290 4922
rect 5314 4870 5344 4922
rect 5344 4870 5356 4922
rect 5356 4870 5370 4922
rect 5394 4870 5408 4922
rect 5408 4870 5420 4922
rect 5420 4870 5450 4922
rect 5474 4870 5484 4922
rect 5484 4870 5530 4922
rect 5234 4868 5290 4870
rect 5314 4868 5370 4870
rect 5394 4868 5450 4870
rect 5474 4868 5530 4870
rect 5234 3834 5290 3836
rect 5314 3834 5370 3836
rect 5394 3834 5450 3836
rect 5474 3834 5530 3836
rect 5234 3782 5280 3834
rect 5280 3782 5290 3834
rect 5314 3782 5344 3834
rect 5344 3782 5356 3834
rect 5356 3782 5370 3834
rect 5394 3782 5408 3834
rect 5408 3782 5420 3834
rect 5420 3782 5450 3834
rect 5474 3782 5484 3834
rect 5484 3782 5530 3834
rect 5234 3780 5290 3782
rect 5314 3780 5370 3782
rect 5394 3780 5450 3782
rect 5474 3780 5530 3782
rect 5998 5616 6054 5652
rect 5894 5466 5950 5468
rect 5974 5466 6030 5468
rect 6054 5466 6110 5468
rect 6134 5466 6190 5468
rect 5894 5414 5940 5466
rect 5940 5414 5950 5466
rect 5974 5414 6004 5466
rect 6004 5414 6016 5466
rect 6016 5414 6030 5466
rect 6054 5414 6068 5466
rect 6068 5414 6080 5466
rect 6080 5414 6110 5466
rect 6134 5414 6144 5466
rect 6144 5414 6190 5466
rect 5894 5412 5950 5414
rect 5974 5412 6030 5414
rect 6054 5412 6110 5414
rect 6134 5412 6190 5414
rect 5894 4378 5950 4380
rect 5974 4378 6030 4380
rect 6054 4378 6110 4380
rect 6134 4378 6190 4380
rect 5894 4326 5940 4378
rect 5940 4326 5950 4378
rect 5974 4326 6004 4378
rect 6004 4326 6016 4378
rect 6016 4326 6030 4378
rect 6054 4326 6068 4378
rect 6068 4326 6080 4378
rect 6080 4326 6110 4378
rect 6134 4326 6144 4378
rect 6144 4326 6190 4378
rect 5894 4324 5950 4326
rect 5974 4324 6030 4326
rect 6054 4324 6110 4326
rect 6134 4324 6190 4326
rect 5894 3290 5950 3292
rect 5974 3290 6030 3292
rect 6054 3290 6110 3292
rect 6134 3290 6190 3292
rect 5894 3238 5940 3290
rect 5940 3238 5950 3290
rect 5974 3238 6004 3290
rect 6004 3238 6016 3290
rect 6016 3238 6030 3290
rect 6054 3238 6068 3290
rect 6068 3238 6080 3290
rect 6080 3238 6110 3290
rect 6134 3238 6144 3290
rect 6144 3238 6190 3290
rect 5894 3236 5950 3238
rect 5974 3236 6030 3238
rect 6054 3236 6110 3238
rect 6134 3236 6190 3238
rect 8482 11056 8538 11092
rect 8086 10362 8142 10364
rect 8166 10362 8222 10364
rect 8246 10362 8302 10364
rect 8326 10362 8382 10364
rect 8086 10310 8132 10362
rect 8132 10310 8142 10362
rect 8166 10310 8196 10362
rect 8196 10310 8208 10362
rect 8208 10310 8222 10362
rect 8246 10310 8260 10362
rect 8260 10310 8272 10362
rect 8272 10310 8302 10362
rect 8326 10310 8336 10362
rect 8336 10310 8382 10362
rect 8086 10308 8142 10310
rect 8166 10308 8222 10310
rect 8246 10308 8302 10310
rect 8326 10308 8382 10310
rect 8086 9274 8142 9276
rect 8166 9274 8222 9276
rect 8246 9274 8302 9276
rect 8326 9274 8382 9276
rect 8086 9222 8132 9274
rect 8132 9222 8142 9274
rect 8166 9222 8196 9274
rect 8196 9222 8208 9274
rect 8208 9222 8222 9274
rect 8246 9222 8260 9274
rect 8260 9222 8272 9274
rect 8272 9222 8302 9274
rect 8326 9222 8336 9274
rect 8336 9222 8382 9274
rect 8086 9220 8142 9222
rect 8166 9220 8222 9222
rect 8246 9220 8302 9222
rect 8326 9220 8382 9222
rect 8746 10906 8802 10908
rect 8826 10906 8882 10908
rect 8906 10906 8962 10908
rect 8986 10906 9042 10908
rect 8746 10854 8792 10906
rect 8792 10854 8802 10906
rect 8826 10854 8856 10906
rect 8856 10854 8868 10906
rect 8868 10854 8882 10906
rect 8906 10854 8920 10906
rect 8920 10854 8932 10906
rect 8932 10854 8962 10906
rect 8986 10854 8996 10906
rect 8996 10854 9042 10906
rect 8746 10852 8802 10854
rect 8826 10852 8882 10854
rect 8906 10852 8962 10854
rect 8986 10852 9042 10854
rect 10938 12538 10994 12540
rect 11018 12538 11074 12540
rect 11098 12538 11154 12540
rect 11178 12538 11234 12540
rect 10938 12486 10984 12538
rect 10984 12486 10994 12538
rect 11018 12486 11048 12538
rect 11048 12486 11060 12538
rect 11060 12486 11074 12538
rect 11098 12486 11112 12538
rect 11112 12486 11124 12538
rect 11124 12486 11154 12538
rect 11178 12486 11188 12538
rect 11188 12486 11234 12538
rect 10938 12484 10994 12486
rect 11018 12484 11074 12486
rect 11098 12484 11154 12486
rect 11178 12484 11234 12486
rect 11598 11994 11654 11996
rect 11678 11994 11734 11996
rect 11758 11994 11814 11996
rect 11838 11994 11894 11996
rect 11598 11942 11644 11994
rect 11644 11942 11654 11994
rect 11678 11942 11708 11994
rect 11708 11942 11720 11994
rect 11720 11942 11734 11994
rect 11758 11942 11772 11994
rect 11772 11942 11784 11994
rect 11784 11942 11814 11994
rect 11838 11942 11848 11994
rect 11848 11942 11894 11994
rect 11598 11940 11654 11942
rect 11678 11940 11734 11942
rect 11758 11940 11814 11942
rect 11838 11940 11894 11942
rect 10938 11450 10994 11452
rect 11018 11450 11074 11452
rect 11098 11450 11154 11452
rect 11178 11450 11234 11452
rect 10938 11398 10984 11450
rect 10984 11398 10994 11450
rect 11018 11398 11048 11450
rect 11048 11398 11060 11450
rect 11060 11398 11074 11450
rect 11098 11398 11112 11450
rect 11112 11398 11124 11450
rect 11124 11398 11154 11450
rect 11178 11398 11188 11450
rect 11188 11398 11234 11450
rect 10938 11396 10994 11398
rect 11018 11396 11074 11398
rect 11098 11396 11154 11398
rect 11178 11396 11234 11398
rect 8746 9818 8802 9820
rect 8826 9818 8882 9820
rect 8906 9818 8962 9820
rect 8986 9818 9042 9820
rect 8746 9766 8792 9818
rect 8792 9766 8802 9818
rect 8826 9766 8856 9818
rect 8856 9766 8868 9818
rect 8868 9766 8882 9818
rect 8906 9766 8920 9818
rect 8920 9766 8932 9818
rect 8932 9766 8962 9818
rect 8986 9766 8996 9818
rect 8996 9766 9042 9818
rect 8746 9764 8802 9766
rect 8826 9764 8882 9766
rect 8906 9764 8962 9766
rect 8986 9764 9042 9766
rect 8086 8186 8142 8188
rect 8166 8186 8222 8188
rect 8246 8186 8302 8188
rect 8326 8186 8382 8188
rect 8086 8134 8132 8186
rect 8132 8134 8142 8186
rect 8166 8134 8196 8186
rect 8196 8134 8208 8186
rect 8208 8134 8222 8186
rect 8246 8134 8260 8186
rect 8260 8134 8272 8186
rect 8272 8134 8302 8186
rect 8326 8134 8336 8186
rect 8336 8134 8382 8186
rect 8086 8132 8142 8134
rect 8166 8132 8222 8134
rect 8246 8132 8302 8134
rect 8326 8132 8382 8134
rect 8086 7098 8142 7100
rect 8166 7098 8222 7100
rect 8246 7098 8302 7100
rect 8326 7098 8382 7100
rect 8086 7046 8132 7098
rect 8132 7046 8142 7098
rect 8166 7046 8196 7098
rect 8196 7046 8208 7098
rect 8208 7046 8222 7098
rect 8246 7046 8260 7098
rect 8260 7046 8272 7098
rect 8272 7046 8302 7098
rect 8326 7046 8336 7098
rect 8336 7046 8382 7098
rect 8086 7044 8142 7046
rect 8166 7044 8222 7046
rect 8246 7044 8302 7046
rect 8326 7044 8382 7046
rect 8086 6010 8142 6012
rect 8166 6010 8222 6012
rect 8246 6010 8302 6012
rect 8326 6010 8382 6012
rect 8086 5958 8132 6010
rect 8132 5958 8142 6010
rect 8166 5958 8196 6010
rect 8196 5958 8208 6010
rect 8208 5958 8222 6010
rect 8246 5958 8260 6010
rect 8260 5958 8272 6010
rect 8272 5958 8302 6010
rect 8326 5958 8336 6010
rect 8336 5958 8382 6010
rect 8086 5956 8142 5958
rect 8166 5956 8222 5958
rect 8246 5956 8302 5958
rect 8326 5956 8382 5958
rect 9770 9424 9826 9480
rect 8746 8730 8802 8732
rect 8826 8730 8882 8732
rect 8906 8730 8962 8732
rect 8986 8730 9042 8732
rect 8746 8678 8792 8730
rect 8792 8678 8802 8730
rect 8826 8678 8856 8730
rect 8856 8678 8868 8730
rect 8868 8678 8882 8730
rect 8906 8678 8920 8730
rect 8920 8678 8932 8730
rect 8932 8678 8962 8730
rect 8986 8678 8996 8730
rect 8996 8678 9042 8730
rect 8746 8676 8802 8678
rect 8826 8676 8882 8678
rect 8906 8676 8962 8678
rect 8986 8676 9042 8678
rect 8746 7642 8802 7644
rect 8826 7642 8882 7644
rect 8906 7642 8962 7644
rect 8986 7642 9042 7644
rect 8746 7590 8792 7642
rect 8792 7590 8802 7642
rect 8826 7590 8856 7642
rect 8856 7590 8868 7642
rect 8868 7590 8882 7642
rect 8906 7590 8920 7642
rect 8920 7590 8932 7642
rect 8932 7590 8962 7642
rect 8986 7590 8996 7642
rect 8996 7590 9042 7642
rect 8746 7588 8802 7590
rect 8826 7588 8882 7590
rect 8906 7588 8962 7590
rect 8986 7588 9042 7590
rect 8746 6554 8802 6556
rect 8826 6554 8882 6556
rect 8906 6554 8962 6556
rect 8986 6554 9042 6556
rect 8746 6502 8792 6554
rect 8792 6502 8802 6554
rect 8826 6502 8856 6554
rect 8856 6502 8868 6554
rect 8868 6502 8882 6554
rect 8906 6502 8920 6554
rect 8920 6502 8932 6554
rect 8932 6502 8962 6554
rect 8986 6502 8996 6554
rect 8996 6502 9042 6554
rect 8746 6500 8802 6502
rect 8826 6500 8882 6502
rect 8906 6500 8962 6502
rect 8986 6500 9042 6502
rect 9862 6160 9918 6216
rect 8746 5466 8802 5468
rect 8826 5466 8882 5468
rect 8906 5466 8962 5468
rect 8986 5466 9042 5468
rect 8746 5414 8792 5466
rect 8792 5414 8802 5466
rect 8826 5414 8856 5466
rect 8856 5414 8868 5466
rect 8868 5414 8882 5466
rect 8906 5414 8920 5466
rect 8920 5414 8932 5466
rect 8932 5414 8962 5466
rect 8986 5414 8996 5466
rect 8996 5414 9042 5466
rect 8746 5412 8802 5414
rect 8826 5412 8882 5414
rect 8906 5412 8962 5414
rect 8986 5412 9042 5414
rect 8086 4922 8142 4924
rect 8166 4922 8222 4924
rect 8246 4922 8302 4924
rect 8326 4922 8382 4924
rect 8086 4870 8132 4922
rect 8132 4870 8142 4922
rect 8166 4870 8196 4922
rect 8196 4870 8208 4922
rect 8208 4870 8222 4922
rect 8246 4870 8260 4922
rect 8260 4870 8272 4922
rect 8272 4870 8302 4922
rect 8326 4870 8336 4922
rect 8336 4870 8382 4922
rect 8086 4868 8142 4870
rect 8166 4868 8222 4870
rect 8246 4868 8302 4870
rect 8326 4868 8382 4870
rect 8746 4378 8802 4380
rect 8826 4378 8882 4380
rect 8906 4378 8962 4380
rect 8986 4378 9042 4380
rect 8746 4326 8792 4378
rect 8792 4326 8802 4378
rect 8826 4326 8856 4378
rect 8856 4326 8868 4378
rect 8868 4326 8882 4378
rect 8906 4326 8920 4378
rect 8920 4326 8932 4378
rect 8932 4326 8962 4378
rect 8986 4326 8996 4378
rect 8996 4326 9042 4378
rect 8746 4324 8802 4326
rect 8826 4324 8882 4326
rect 8906 4324 8962 4326
rect 8986 4324 9042 4326
rect 8086 3834 8142 3836
rect 8166 3834 8222 3836
rect 8246 3834 8302 3836
rect 8326 3834 8382 3836
rect 8086 3782 8132 3834
rect 8132 3782 8142 3834
rect 8166 3782 8196 3834
rect 8196 3782 8208 3834
rect 8208 3782 8222 3834
rect 8246 3782 8260 3834
rect 8260 3782 8272 3834
rect 8272 3782 8302 3834
rect 8326 3782 8336 3834
rect 8336 3782 8382 3834
rect 8086 3780 8142 3782
rect 8166 3780 8222 3782
rect 8246 3780 8302 3782
rect 8326 3780 8382 3782
rect 5234 2746 5290 2748
rect 5314 2746 5370 2748
rect 5394 2746 5450 2748
rect 5474 2746 5530 2748
rect 5234 2694 5280 2746
rect 5280 2694 5290 2746
rect 5314 2694 5344 2746
rect 5344 2694 5356 2746
rect 5356 2694 5370 2746
rect 5394 2694 5408 2746
rect 5408 2694 5420 2746
rect 5420 2694 5450 2746
rect 5474 2694 5484 2746
rect 5484 2694 5530 2746
rect 5234 2692 5290 2694
rect 5314 2692 5370 2694
rect 5394 2692 5450 2694
rect 5474 2692 5530 2694
rect 3042 2202 3098 2204
rect 3122 2202 3178 2204
rect 3202 2202 3258 2204
rect 3282 2202 3338 2204
rect 3042 2150 3088 2202
rect 3088 2150 3098 2202
rect 3122 2150 3152 2202
rect 3152 2150 3164 2202
rect 3164 2150 3178 2202
rect 3202 2150 3216 2202
rect 3216 2150 3228 2202
rect 3228 2150 3258 2202
rect 3282 2150 3292 2202
rect 3292 2150 3338 2202
rect 3042 2148 3098 2150
rect 3122 2148 3178 2150
rect 3202 2148 3258 2150
rect 3282 2148 3338 2150
rect 8086 2746 8142 2748
rect 8166 2746 8222 2748
rect 8246 2746 8302 2748
rect 8326 2746 8382 2748
rect 8086 2694 8132 2746
rect 8132 2694 8142 2746
rect 8166 2694 8196 2746
rect 8196 2694 8208 2746
rect 8208 2694 8222 2746
rect 8246 2694 8260 2746
rect 8260 2694 8272 2746
rect 8272 2694 8302 2746
rect 8326 2694 8336 2746
rect 8336 2694 8382 2746
rect 8086 2692 8142 2694
rect 8166 2692 8222 2694
rect 8246 2692 8302 2694
rect 8326 2692 8382 2694
rect 8746 3290 8802 3292
rect 8826 3290 8882 3292
rect 8906 3290 8962 3292
rect 8986 3290 9042 3292
rect 8746 3238 8792 3290
rect 8792 3238 8802 3290
rect 8826 3238 8856 3290
rect 8856 3238 8868 3290
rect 8868 3238 8882 3290
rect 8906 3238 8920 3290
rect 8920 3238 8932 3290
rect 8932 3238 8962 3290
rect 8986 3238 8996 3290
rect 8996 3238 9042 3290
rect 8746 3236 8802 3238
rect 8826 3236 8882 3238
rect 8906 3236 8962 3238
rect 8986 3236 9042 3238
rect 11598 10906 11654 10908
rect 11678 10906 11734 10908
rect 11758 10906 11814 10908
rect 11838 10906 11894 10908
rect 11598 10854 11644 10906
rect 11644 10854 11654 10906
rect 11678 10854 11708 10906
rect 11708 10854 11720 10906
rect 11720 10854 11734 10906
rect 11758 10854 11772 10906
rect 11772 10854 11784 10906
rect 11784 10854 11814 10906
rect 11838 10854 11848 10906
rect 11848 10854 11894 10906
rect 11598 10852 11654 10854
rect 11678 10852 11734 10854
rect 11758 10852 11814 10854
rect 11838 10852 11894 10854
rect 10938 10362 10994 10364
rect 11018 10362 11074 10364
rect 11098 10362 11154 10364
rect 11178 10362 11234 10364
rect 10938 10310 10984 10362
rect 10984 10310 10994 10362
rect 11018 10310 11048 10362
rect 11048 10310 11060 10362
rect 11060 10310 11074 10362
rect 11098 10310 11112 10362
rect 11112 10310 11124 10362
rect 11124 10310 11154 10362
rect 11178 10310 11188 10362
rect 11188 10310 11234 10362
rect 10938 10308 10994 10310
rect 11018 10308 11074 10310
rect 11098 10308 11154 10310
rect 11178 10308 11234 10310
rect 10938 9274 10994 9276
rect 11018 9274 11074 9276
rect 11098 9274 11154 9276
rect 11178 9274 11234 9276
rect 10938 9222 10984 9274
rect 10984 9222 10994 9274
rect 11018 9222 11048 9274
rect 11048 9222 11060 9274
rect 11060 9222 11074 9274
rect 11098 9222 11112 9274
rect 11112 9222 11124 9274
rect 11124 9222 11154 9274
rect 11178 9222 11188 9274
rect 11188 9222 11234 9274
rect 10938 9220 10994 9222
rect 11018 9220 11074 9222
rect 11098 9220 11154 9222
rect 11178 9220 11234 9222
rect 10938 8186 10994 8188
rect 11018 8186 11074 8188
rect 11098 8186 11154 8188
rect 11178 8186 11234 8188
rect 10938 8134 10984 8186
rect 10984 8134 10994 8186
rect 11018 8134 11048 8186
rect 11048 8134 11060 8186
rect 11060 8134 11074 8186
rect 11098 8134 11112 8186
rect 11112 8134 11124 8186
rect 11124 8134 11154 8186
rect 11178 8134 11188 8186
rect 11188 8134 11234 8186
rect 10938 8132 10994 8134
rect 11018 8132 11074 8134
rect 11098 8132 11154 8134
rect 11178 8132 11234 8134
rect 11598 9818 11654 9820
rect 11678 9818 11734 9820
rect 11758 9818 11814 9820
rect 11838 9818 11894 9820
rect 11598 9766 11644 9818
rect 11644 9766 11654 9818
rect 11678 9766 11708 9818
rect 11708 9766 11720 9818
rect 11720 9766 11734 9818
rect 11758 9766 11772 9818
rect 11772 9766 11784 9818
rect 11784 9766 11814 9818
rect 11838 9766 11848 9818
rect 11848 9766 11894 9818
rect 11598 9764 11654 9766
rect 11678 9764 11734 9766
rect 11758 9764 11814 9766
rect 11838 9764 11894 9766
rect 11598 8730 11654 8732
rect 11678 8730 11734 8732
rect 11758 8730 11814 8732
rect 11838 8730 11894 8732
rect 11598 8678 11644 8730
rect 11644 8678 11654 8730
rect 11678 8678 11708 8730
rect 11708 8678 11720 8730
rect 11720 8678 11734 8730
rect 11758 8678 11772 8730
rect 11772 8678 11784 8730
rect 11784 8678 11814 8730
rect 11838 8678 11848 8730
rect 11848 8678 11894 8730
rect 11598 8676 11654 8678
rect 11678 8676 11734 8678
rect 11758 8676 11814 8678
rect 11838 8676 11894 8678
rect 11598 7642 11654 7644
rect 11678 7642 11734 7644
rect 11758 7642 11814 7644
rect 11838 7642 11894 7644
rect 11598 7590 11644 7642
rect 11644 7590 11654 7642
rect 11678 7590 11708 7642
rect 11708 7590 11720 7642
rect 11720 7590 11734 7642
rect 11758 7590 11772 7642
rect 11772 7590 11784 7642
rect 11784 7590 11814 7642
rect 11838 7590 11848 7642
rect 11848 7590 11894 7642
rect 11598 7588 11654 7590
rect 11678 7588 11734 7590
rect 11758 7588 11814 7590
rect 11838 7588 11894 7590
rect 12070 8880 12126 8936
rect 10938 7098 10994 7100
rect 11018 7098 11074 7100
rect 11098 7098 11154 7100
rect 11178 7098 11234 7100
rect 10938 7046 10984 7098
rect 10984 7046 10994 7098
rect 11018 7046 11048 7098
rect 11048 7046 11060 7098
rect 11060 7046 11074 7098
rect 11098 7046 11112 7098
rect 11112 7046 11124 7098
rect 11124 7046 11154 7098
rect 11178 7046 11188 7098
rect 11188 7046 11234 7098
rect 10938 7044 10994 7046
rect 11018 7044 11074 7046
rect 11098 7044 11154 7046
rect 11178 7044 11234 7046
rect 11598 6554 11654 6556
rect 11678 6554 11734 6556
rect 11758 6554 11814 6556
rect 11838 6554 11894 6556
rect 11598 6502 11644 6554
rect 11644 6502 11654 6554
rect 11678 6502 11708 6554
rect 11708 6502 11720 6554
rect 11720 6502 11734 6554
rect 11758 6502 11772 6554
rect 11772 6502 11784 6554
rect 11784 6502 11814 6554
rect 11838 6502 11848 6554
rect 11848 6502 11894 6554
rect 11598 6500 11654 6502
rect 11678 6500 11734 6502
rect 11758 6500 11814 6502
rect 11838 6500 11894 6502
rect 12162 6860 12218 6896
rect 12162 6840 12164 6860
rect 12164 6840 12216 6860
rect 12216 6840 12218 6860
rect 11610 6180 11666 6216
rect 11610 6160 11612 6180
rect 11612 6160 11664 6180
rect 11664 6160 11666 6180
rect 10938 6010 10994 6012
rect 11018 6010 11074 6012
rect 11098 6010 11154 6012
rect 11178 6010 11234 6012
rect 10938 5958 10984 6010
rect 10984 5958 10994 6010
rect 11018 5958 11048 6010
rect 11048 5958 11060 6010
rect 11060 5958 11074 6010
rect 11098 5958 11112 6010
rect 11112 5958 11124 6010
rect 11124 5958 11154 6010
rect 11178 5958 11188 6010
rect 11188 5958 11234 6010
rect 10938 5956 10994 5958
rect 11018 5956 11074 5958
rect 11098 5956 11154 5958
rect 11178 5956 11234 5958
rect 11598 5466 11654 5468
rect 11678 5466 11734 5468
rect 11758 5466 11814 5468
rect 11838 5466 11894 5468
rect 11598 5414 11644 5466
rect 11644 5414 11654 5466
rect 11678 5414 11708 5466
rect 11708 5414 11720 5466
rect 11720 5414 11734 5466
rect 11758 5414 11772 5466
rect 11772 5414 11784 5466
rect 11784 5414 11814 5466
rect 11838 5414 11848 5466
rect 11848 5414 11894 5466
rect 11598 5412 11654 5414
rect 11678 5412 11734 5414
rect 11758 5412 11814 5414
rect 11838 5412 11894 5414
rect 10938 4922 10994 4924
rect 11018 4922 11074 4924
rect 11098 4922 11154 4924
rect 11178 4922 11234 4924
rect 10938 4870 10984 4922
rect 10984 4870 10994 4922
rect 11018 4870 11048 4922
rect 11048 4870 11060 4922
rect 11060 4870 11074 4922
rect 11098 4870 11112 4922
rect 11112 4870 11124 4922
rect 11124 4870 11154 4922
rect 11178 4870 11188 4922
rect 11188 4870 11234 4922
rect 10938 4868 10994 4870
rect 11018 4868 11074 4870
rect 11098 4868 11154 4870
rect 11178 4868 11234 4870
rect 11702 4800 11758 4856
rect 12070 6160 12126 6216
rect 12162 5480 12218 5536
rect 11598 4378 11654 4380
rect 11678 4378 11734 4380
rect 11758 4378 11814 4380
rect 11838 4378 11894 4380
rect 11598 4326 11644 4378
rect 11644 4326 11654 4378
rect 11678 4326 11708 4378
rect 11708 4326 11720 4378
rect 11720 4326 11734 4378
rect 11758 4326 11772 4378
rect 11772 4326 11784 4378
rect 11784 4326 11814 4378
rect 11838 4326 11848 4378
rect 11848 4326 11894 4378
rect 11598 4324 11654 4326
rect 11678 4324 11734 4326
rect 11758 4324 11814 4326
rect 11838 4324 11894 4326
rect 10938 3834 10994 3836
rect 11018 3834 11074 3836
rect 11098 3834 11154 3836
rect 11178 3834 11234 3836
rect 10938 3782 10984 3834
rect 10984 3782 10994 3834
rect 11018 3782 11048 3834
rect 11048 3782 11060 3834
rect 11060 3782 11074 3834
rect 11098 3782 11112 3834
rect 11112 3782 11124 3834
rect 11124 3782 11154 3834
rect 11178 3782 11188 3834
rect 11188 3782 11234 3834
rect 10938 3780 10994 3782
rect 11018 3780 11074 3782
rect 11098 3780 11154 3782
rect 11178 3780 11234 3782
rect 11598 3290 11654 3292
rect 11678 3290 11734 3292
rect 11758 3290 11814 3292
rect 11838 3290 11894 3292
rect 11598 3238 11644 3290
rect 11644 3238 11654 3290
rect 11678 3238 11708 3290
rect 11708 3238 11720 3290
rect 11720 3238 11734 3290
rect 11758 3238 11772 3290
rect 11772 3238 11784 3290
rect 11784 3238 11814 3290
rect 11838 3238 11848 3290
rect 11848 3238 11894 3290
rect 11598 3236 11654 3238
rect 11678 3236 11734 3238
rect 11758 3236 11814 3238
rect 11838 3236 11894 3238
rect 10938 2746 10994 2748
rect 11018 2746 11074 2748
rect 11098 2746 11154 2748
rect 11178 2746 11234 2748
rect 10938 2694 10984 2746
rect 10984 2694 10994 2746
rect 11018 2694 11048 2746
rect 11048 2694 11060 2746
rect 11060 2694 11074 2746
rect 11098 2694 11112 2746
rect 11112 2694 11124 2746
rect 11124 2694 11154 2746
rect 11178 2694 11188 2746
rect 11188 2694 11234 2746
rect 10938 2692 10994 2694
rect 11018 2692 11074 2694
rect 11098 2692 11154 2694
rect 11178 2692 11234 2694
rect 5894 2202 5950 2204
rect 5974 2202 6030 2204
rect 6054 2202 6110 2204
rect 6134 2202 6190 2204
rect 5894 2150 5940 2202
rect 5940 2150 5950 2202
rect 5974 2150 6004 2202
rect 6004 2150 6016 2202
rect 6016 2150 6030 2202
rect 6054 2150 6068 2202
rect 6068 2150 6080 2202
rect 6080 2150 6110 2202
rect 6134 2150 6144 2202
rect 6144 2150 6190 2202
rect 5894 2148 5950 2150
rect 5974 2148 6030 2150
rect 6054 2148 6110 2150
rect 6134 2148 6190 2150
rect 8746 2202 8802 2204
rect 8826 2202 8882 2204
rect 8906 2202 8962 2204
rect 8986 2202 9042 2204
rect 8746 2150 8792 2202
rect 8792 2150 8802 2202
rect 8826 2150 8856 2202
rect 8856 2150 8868 2202
rect 8868 2150 8882 2202
rect 8906 2150 8920 2202
rect 8920 2150 8932 2202
rect 8932 2150 8962 2202
rect 8986 2150 8996 2202
rect 8996 2150 9042 2202
rect 8746 2148 8802 2150
rect 8826 2148 8882 2150
rect 8906 2148 8962 2150
rect 8986 2148 9042 2150
rect 11598 2202 11654 2204
rect 11678 2202 11734 2204
rect 11758 2202 11814 2204
rect 11838 2202 11894 2204
rect 11598 2150 11644 2202
rect 11644 2150 11654 2202
rect 11678 2150 11708 2202
rect 11708 2150 11720 2202
rect 11720 2150 11734 2202
rect 11758 2150 11772 2202
rect 11772 2150 11784 2202
rect 11784 2150 11814 2202
rect 11838 2150 11848 2202
rect 11848 2150 11894 2202
rect 11598 2148 11654 2150
rect 11678 2148 11734 2150
rect 11758 2148 11814 2150
rect 11838 2148 11894 2150
<< metal3 >>
rect 2372 13632 2688 13633
rect 2372 13568 2378 13632
rect 2442 13568 2458 13632
rect 2522 13568 2538 13632
rect 2602 13568 2618 13632
rect 2682 13568 2688 13632
rect 2372 13567 2688 13568
rect 5224 13632 5540 13633
rect 5224 13568 5230 13632
rect 5294 13568 5310 13632
rect 5374 13568 5390 13632
rect 5454 13568 5470 13632
rect 5534 13568 5540 13632
rect 5224 13567 5540 13568
rect 8076 13632 8392 13633
rect 8076 13568 8082 13632
rect 8146 13568 8162 13632
rect 8226 13568 8242 13632
rect 8306 13568 8322 13632
rect 8386 13568 8392 13632
rect 8076 13567 8392 13568
rect 10928 13632 11244 13633
rect 10928 13568 10934 13632
rect 10998 13568 11014 13632
rect 11078 13568 11094 13632
rect 11158 13568 11174 13632
rect 11238 13568 11244 13632
rect 10928 13567 11244 13568
rect 3032 13088 3348 13089
rect 3032 13024 3038 13088
rect 3102 13024 3118 13088
rect 3182 13024 3198 13088
rect 3262 13024 3278 13088
rect 3342 13024 3348 13088
rect 3032 13023 3348 13024
rect 5884 13088 6200 13089
rect 5884 13024 5890 13088
rect 5954 13024 5970 13088
rect 6034 13024 6050 13088
rect 6114 13024 6130 13088
rect 6194 13024 6200 13088
rect 5884 13023 6200 13024
rect 8736 13088 9052 13089
rect 8736 13024 8742 13088
rect 8806 13024 8822 13088
rect 8886 13024 8902 13088
rect 8966 13024 8982 13088
rect 9046 13024 9052 13088
rect 8736 13023 9052 13024
rect 11588 13088 11904 13089
rect 11588 13024 11594 13088
rect 11658 13024 11674 13088
rect 11738 13024 11754 13088
rect 11818 13024 11834 13088
rect 11898 13024 11904 13088
rect 11588 13023 11904 13024
rect 2372 12544 2688 12545
rect 2372 12480 2378 12544
rect 2442 12480 2458 12544
rect 2522 12480 2538 12544
rect 2602 12480 2618 12544
rect 2682 12480 2688 12544
rect 2372 12479 2688 12480
rect 5224 12544 5540 12545
rect 5224 12480 5230 12544
rect 5294 12480 5310 12544
rect 5374 12480 5390 12544
rect 5454 12480 5470 12544
rect 5534 12480 5540 12544
rect 5224 12479 5540 12480
rect 8076 12544 8392 12545
rect 8076 12480 8082 12544
rect 8146 12480 8162 12544
rect 8226 12480 8242 12544
rect 8306 12480 8322 12544
rect 8386 12480 8392 12544
rect 8076 12479 8392 12480
rect 10928 12544 11244 12545
rect 10928 12480 10934 12544
rect 10998 12480 11014 12544
rect 11078 12480 11094 12544
rect 11158 12480 11174 12544
rect 11238 12480 11244 12544
rect 10928 12479 11244 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 4521 12202 4587 12205
rect 5257 12202 5323 12205
rect 4521 12200 5323 12202
rect 4521 12144 4526 12200
rect 4582 12144 5262 12200
rect 5318 12144 5323 12200
rect 4521 12142 5323 12144
rect 4521 12139 4587 12142
rect 5257 12139 5323 12142
rect 3032 12000 3348 12001
rect 3032 11936 3038 12000
rect 3102 11936 3118 12000
rect 3182 11936 3198 12000
rect 3262 11936 3278 12000
rect 3342 11936 3348 12000
rect 3032 11935 3348 11936
rect 5884 12000 6200 12001
rect 5884 11936 5890 12000
rect 5954 11936 5970 12000
rect 6034 11936 6050 12000
rect 6114 11936 6130 12000
rect 6194 11936 6200 12000
rect 5884 11935 6200 11936
rect 8736 12000 9052 12001
rect 8736 11936 8742 12000
rect 8806 11936 8822 12000
rect 8886 11936 8902 12000
rect 8966 11936 8982 12000
rect 9046 11936 9052 12000
rect 8736 11935 9052 11936
rect 11588 12000 11904 12001
rect 11588 11936 11594 12000
rect 11658 11936 11674 12000
rect 11738 11936 11754 12000
rect 11818 11936 11834 12000
rect 11898 11936 11904 12000
rect 11588 11935 11904 11936
rect 0 11658 800 11688
rect 1025 11658 1091 11661
rect 0 11656 1091 11658
rect 0 11600 1030 11656
rect 1086 11600 1091 11656
rect 0 11598 1091 11600
rect 0 11568 800 11598
rect 1025 11595 1091 11598
rect 2372 11456 2688 11457
rect 2372 11392 2378 11456
rect 2442 11392 2458 11456
rect 2522 11392 2538 11456
rect 2602 11392 2618 11456
rect 2682 11392 2688 11456
rect 2372 11391 2688 11392
rect 5224 11456 5540 11457
rect 5224 11392 5230 11456
rect 5294 11392 5310 11456
rect 5374 11392 5390 11456
rect 5454 11392 5470 11456
rect 5534 11392 5540 11456
rect 5224 11391 5540 11392
rect 8076 11456 8392 11457
rect 8076 11392 8082 11456
rect 8146 11392 8162 11456
rect 8226 11392 8242 11456
rect 8306 11392 8322 11456
rect 8386 11392 8392 11456
rect 8076 11391 8392 11392
rect 10928 11456 11244 11457
rect 10928 11392 10934 11456
rect 10998 11392 11014 11456
rect 11078 11392 11094 11456
rect 11158 11392 11174 11456
rect 11238 11392 11244 11456
rect 10928 11391 11244 11392
rect 7649 11114 7715 11117
rect 8477 11114 8543 11117
rect 7649 11112 8543 11114
rect 7649 11056 7654 11112
rect 7710 11056 8482 11112
rect 8538 11056 8543 11112
rect 7649 11054 8543 11056
rect 7649 11051 7715 11054
rect 8477 11051 8543 11054
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 3032 10912 3348 10913
rect 3032 10848 3038 10912
rect 3102 10848 3118 10912
rect 3182 10848 3198 10912
rect 3262 10848 3278 10912
rect 3342 10848 3348 10912
rect 3032 10847 3348 10848
rect 5884 10912 6200 10913
rect 5884 10848 5890 10912
rect 5954 10848 5970 10912
rect 6034 10848 6050 10912
rect 6114 10848 6130 10912
rect 6194 10848 6200 10912
rect 5884 10847 6200 10848
rect 8736 10912 9052 10913
rect 8736 10848 8742 10912
rect 8806 10848 8822 10912
rect 8886 10848 8902 10912
rect 8966 10848 8982 10912
rect 9046 10848 9052 10912
rect 8736 10847 9052 10848
rect 11588 10912 11904 10913
rect 11588 10848 11594 10912
rect 11658 10848 11674 10912
rect 11738 10848 11754 10912
rect 11818 10848 11834 10912
rect 11898 10848 11904 10912
rect 11588 10847 11904 10848
rect 2372 10368 2688 10369
rect 2372 10304 2378 10368
rect 2442 10304 2458 10368
rect 2522 10304 2538 10368
rect 2602 10304 2618 10368
rect 2682 10304 2688 10368
rect 2372 10303 2688 10304
rect 5224 10368 5540 10369
rect 5224 10304 5230 10368
rect 5294 10304 5310 10368
rect 5374 10304 5390 10368
rect 5454 10304 5470 10368
rect 5534 10304 5540 10368
rect 5224 10303 5540 10304
rect 8076 10368 8392 10369
rect 8076 10304 8082 10368
rect 8146 10304 8162 10368
rect 8226 10304 8242 10368
rect 8306 10304 8322 10368
rect 8386 10304 8392 10368
rect 8076 10303 8392 10304
rect 10928 10368 11244 10369
rect 10928 10304 10934 10368
rect 10998 10304 11014 10368
rect 11078 10304 11094 10368
rect 11158 10304 11174 10368
rect 11238 10304 11244 10368
rect 10928 10303 11244 10304
rect 3032 9824 3348 9825
rect 3032 9760 3038 9824
rect 3102 9760 3118 9824
rect 3182 9760 3198 9824
rect 3262 9760 3278 9824
rect 3342 9760 3348 9824
rect 3032 9759 3348 9760
rect 5884 9824 6200 9825
rect 5884 9760 5890 9824
rect 5954 9760 5970 9824
rect 6034 9760 6050 9824
rect 6114 9760 6130 9824
rect 6194 9760 6200 9824
rect 5884 9759 6200 9760
rect 8736 9824 9052 9825
rect 8736 9760 8742 9824
rect 8806 9760 8822 9824
rect 8886 9760 8902 9824
rect 8966 9760 8982 9824
rect 9046 9760 9052 9824
rect 8736 9759 9052 9760
rect 11588 9824 11904 9825
rect 11588 9760 11594 9824
rect 11658 9760 11674 9824
rect 11738 9760 11754 9824
rect 11818 9760 11834 9824
rect 11898 9760 11904 9824
rect 11588 9759 11904 9760
rect 1669 9618 1735 9621
rect 3141 9618 3207 9621
rect 1669 9616 3207 9618
rect 1669 9560 1674 9616
rect 1730 9560 3146 9616
rect 3202 9560 3207 9616
rect 1669 9558 3207 9560
rect 1669 9555 1735 9558
rect 3141 9555 3207 9558
rect 2589 9482 2655 9485
rect 9765 9482 9831 9485
rect 2589 9480 9831 9482
rect 2589 9424 2594 9480
rect 2650 9424 9770 9480
rect 9826 9424 9831 9480
rect 2589 9422 9831 9424
rect 2589 9419 2655 9422
rect 9765 9419 9831 9422
rect 2372 9280 2688 9281
rect 2372 9216 2378 9280
rect 2442 9216 2458 9280
rect 2522 9216 2538 9280
rect 2602 9216 2618 9280
rect 2682 9216 2688 9280
rect 2372 9215 2688 9216
rect 5224 9280 5540 9281
rect 5224 9216 5230 9280
rect 5294 9216 5310 9280
rect 5374 9216 5390 9280
rect 5454 9216 5470 9280
rect 5534 9216 5540 9280
rect 5224 9215 5540 9216
rect 8076 9280 8392 9281
rect 8076 9216 8082 9280
rect 8146 9216 8162 9280
rect 8226 9216 8242 9280
rect 8306 9216 8322 9280
rect 8386 9216 8392 9280
rect 8076 9215 8392 9216
rect 10928 9280 11244 9281
rect 10928 9216 10934 9280
rect 10998 9216 11014 9280
rect 11078 9216 11094 9280
rect 11158 9216 11174 9280
rect 11238 9216 11244 9280
rect 10928 9215 11244 9216
rect 1485 9074 1551 9077
rect 2221 9074 2287 9077
rect 4245 9074 4311 9077
rect 1485 9072 4311 9074
rect 1485 9016 1490 9072
rect 1546 9016 2226 9072
rect 2282 9016 4250 9072
rect 4306 9016 4311 9072
rect 1485 9014 4311 9016
rect 1485 9011 1551 9014
rect 2221 9011 2287 9014
rect 4245 9011 4311 9014
rect 0 8938 800 8968
rect 1485 8938 1551 8941
rect 0 8936 1551 8938
rect 0 8880 1490 8936
rect 1546 8880 1551 8936
rect 0 8878 1551 8880
rect 0 8848 800 8878
rect 1485 8875 1551 8878
rect 12065 8938 12131 8941
rect 12846 8938 13646 8968
rect 12065 8936 13646 8938
rect 12065 8880 12070 8936
rect 12126 8880 13646 8936
rect 12065 8878 13646 8880
rect 12065 8875 12131 8878
rect 12846 8848 13646 8878
rect 3032 8736 3348 8737
rect 3032 8672 3038 8736
rect 3102 8672 3118 8736
rect 3182 8672 3198 8736
rect 3262 8672 3278 8736
rect 3342 8672 3348 8736
rect 3032 8671 3348 8672
rect 5884 8736 6200 8737
rect 5884 8672 5890 8736
rect 5954 8672 5970 8736
rect 6034 8672 6050 8736
rect 6114 8672 6130 8736
rect 6194 8672 6200 8736
rect 5884 8671 6200 8672
rect 8736 8736 9052 8737
rect 8736 8672 8742 8736
rect 8806 8672 8822 8736
rect 8886 8672 8902 8736
rect 8966 8672 8982 8736
rect 9046 8672 9052 8736
rect 8736 8671 9052 8672
rect 11588 8736 11904 8737
rect 11588 8672 11594 8736
rect 11658 8672 11674 8736
rect 11738 8672 11754 8736
rect 11818 8672 11834 8736
rect 11898 8672 11904 8736
rect 11588 8671 11904 8672
rect 2589 8530 2655 8533
rect 4889 8530 4955 8533
rect 2589 8528 4955 8530
rect 2589 8472 2594 8528
rect 2650 8472 4894 8528
rect 4950 8472 4955 8528
rect 2589 8470 4955 8472
rect 2589 8467 2655 8470
rect 4889 8467 4955 8470
rect 3141 8394 3207 8397
rect 4521 8394 4587 8397
rect 3141 8392 4587 8394
rect 3141 8336 3146 8392
rect 3202 8336 4526 8392
rect 4582 8336 4587 8392
rect 3141 8334 4587 8336
rect 3141 8331 3207 8334
rect 4521 8331 4587 8334
rect 0 8258 800 8288
rect 1301 8258 1367 8261
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 0 8168 800 8198
rect 1301 8195 1367 8198
rect 2372 8192 2688 8193
rect 2372 8128 2378 8192
rect 2442 8128 2458 8192
rect 2522 8128 2538 8192
rect 2602 8128 2618 8192
rect 2682 8128 2688 8192
rect 2372 8127 2688 8128
rect 5224 8192 5540 8193
rect 5224 8128 5230 8192
rect 5294 8128 5310 8192
rect 5374 8128 5390 8192
rect 5454 8128 5470 8192
rect 5534 8128 5540 8192
rect 5224 8127 5540 8128
rect 8076 8192 8392 8193
rect 8076 8128 8082 8192
rect 8146 8128 8162 8192
rect 8226 8128 8242 8192
rect 8306 8128 8322 8192
rect 8386 8128 8392 8192
rect 8076 8127 8392 8128
rect 10928 8192 11244 8193
rect 10928 8128 10934 8192
rect 10998 8128 11014 8192
rect 11078 8128 11094 8192
rect 11158 8128 11174 8192
rect 11238 8128 11244 8192
rect 10928 8127 11244 8128
rect 3032 7648 3348 7649
rect 0 7578 800 7608
rect 3032 7584 3038 7648
rect 3102 7584 3118 7648
rect 3182 7584 3198 7648
rect 3262 7584 3278 7648
rect 3342 7584 3348 7648
rect 3032 7583 3348 7584
rect 5884 7648 6200 7649
rect 5884 7584 5890 7648
rect 5954 7584 5970 7648
rect 6034 7584 6050 7648
rect 6114 7584 6130 7648
rect 6194 7584 6200 7648
rect 5884 7583 6200 7584
rect 8736 7648 9052 7649
rect 8736 7584 8742 7648
rect 8806 7584 8822 7648
rect 8886 7584 8902 7648
rect 8966 7584 8982 7648
rect 9046 7584 9052 7648
rect 8736 7583 9052 7584
rect 11588 7648 11904 7649
rect 11588 7584 11594 7648
rect 11658 7584 11674 7648
rect 11738 7584 11754 7648
rect 11818 7584 11834 7648
rect 11898 7584 11904 7648
rect 11588 7583 11904 7584
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 2372 7104 2688 7105
rect 2372 7040 2378 7104
rect 2442 7040 2458 7104
rect 2522 7040 2538 7104
rect 2602 7040 2618 7104
rect 2682 7040 2688 7104
rect 2372 7039 2688 7040
rect 5224 7104 5540 7105
rect 5224 7040 5230 7104
rect 5294 7040 5310 7104
rect 5374 7040 5390 7104
rect 5454 7040 5470 7104
rect 5534 7040 5540 7104
rect 5224 7039 5540 7040
rect 8076 7104 8392 7105
rect 8076 7040 8082 7104
rect 8146 7040 8162 7104
rect 8226 7040 8242 7104
rect 8306 7040 8322 7104
rect 8386 7040 8392 7104
rect 8076 7039 8392 7040
rect 10928 7104 11244 7105
rect 10928 7040 10934 7104
rect 10998 7040 11014 7104
rect 11078 7040 11094 7104
rect 11158 7040 11174 7104
rect 11238 7040 11244 7104
rect 10928 7039 11244 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 12157 6898 12223 6901
rect 12846 6898 13646 6928
rect 12157 6896 13646 6898
rect 12157 6840 12162 6896
rect 12218 6840 13646 6896
rect 12157 6838 13646 6840
rect 12157 6835 12223 6838
rect 12846 6808 13646 6838
rect 3032 6560 3348 6561
rect 3032 6496 3038 6560
rect 3102 6496 3118 6560
rect 3182 6496 3198 6560
rect 3262 6496 3278 6560
rect 3342 6496 3348 6560
rect 3032 6495 3348 6496
rect 5884 6560 6200 6561
rect 5884 6496 5890 6560
rect 5954 6496 5970 6560
rect 6034 6496 6050 6560
rect 6114 6496 6130 6560
rect 6194 6496 6200 6560
rect 5884 6495 6200 6496
rect 8736 6560 9052 6561
rect 8736 6496 8742 6560
rect 8806 6496 8822 6560
rect 8886 6496 8902 6560
rect 8966 6496 8982 6560
rect 9046 6496 9052 6560
rect 8736 6495 9052 6496
rect 11588 6560 11904 6561
rect 11588 6496 11594 6560
rect 11658 6496 11674 6560
rect 11738 6496 11754 6560
rect 11818 6496 11834 6560
rect 11898 6496 11904 6560
rect 11588 6495 11904 6496
rect 0 6218 800 6248
rect 9857 6218 9923 6221
rect 11605 6218 11671 6221
rect 0 6128 858 6218
rect 9857 6216 11671 6218
rect 9857 6160 9862 6216
rect 9918 6160 11610 6216
rect 11666 6160 11671 6216
rect 9857 6158 11671 6160
rect 9857 6155 9923 6158
rect 11605 6155 11671 6158
rect 12065 6218 12131 6221
rect 12846 6218 13646 6248
rect 12065 6216 13646 6218
rect 12065 6160 12070 6216
rect 12126 6160 13646 6216
rect 12065 6158 13646 6160
rect 12065 6155 12131 6158
rect 12846 6128 13646 6158
rect 798 6085 858 6128
rect 798 6080 907 6085
rect 798 6024 846 6080
rect 902 6024 907 6080
rect 798 6022 907 6024
rect 841 6019 907 6022
rect 2372 6016 2688 6017
rect 2372 5952 2378 6016
rect 2442 5952 2458 6016
rect 2522 5952 2538 6016
rect 2602 5952 2618 6016
rect 2682 5952 2688 6016
rect 2372 5951 2688 5952
rect 5224 6016 5540 6017
rect 5224 5952 5230 6016
rect 5294 5952 5310 6016
rect 5374 5952 5390 6016
rect 5454 5952 5470 6016
rect 5534 5952 5540 6016
rect 5224 5951 5540 5952
rect 8076 6016 8392 6017
rect 8076 5952 8082 6016
rect 8146 5952 8162 6016
rect 8226 5952 8242 6016
rect 8306 5952 8322 6016
rect 8386 5952 8392 6016
rect 8076 5951 8392 5952
rect 10928 6016 11244 6017
rect 10928 5952 10934 6016
rect 10998 5952 11014 6016
rect 11078 5952 11094 6016
rect 11158 5952 11174 6016
rect 11238 5952 11244 6016
rect 10928 5951 11244 5952
rect 4153 5674 4219 5677
rect 5993 5674 6059 5677
rect 4153 5672 6059 5674
rect 4153 5616 4158 5672
rect 4214 5616 5998 5672
rect 6054 5616 6059 5672
rect 4153 5614 6059 5616
rect 4153 5611 4219 5614
rect 5993 5611 6059 5614
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 12157 5538 12223 5541
rect 12846 5538 13646 5568
rect 12157 5536 13646 5538
rect 12157 5480 12162 5536
rect 12218 5480 13646 5536
rect 12157 5478 13646 5480
rect 12157 5475 12223 5478
rect 3032 5472 3348 5473
rect 3032 5408 3038 5472
rect 3102 5408 3118 5472
rect 3182 5408 3198 5472
rect 3262 5408 3278 5472
rect 3342 5408 3348 5472
rect 3032 5407 3348 5408
rect 5884 5472 6200 5473
rect 5884 5408 5890 5472
rect 5954 5408 5970 5472
rect 6034 5408 6050 5472
rect 6114 5408 6130 5472
rect 6194 5408 6200 5472
rect 5884 5407 6200 5408
rect 8736 5472 9052 5473
rect 8736 5408 8742 5472
rect 8806 5408 8822 5472
rect 8886 5408 8902 5472
rect 8966 5408 8982 5472
rect 9046 5408 9052 5472
rect 8736 5407 9052 5408
rect 11588 5472 11904 5473
rect 11588 5408 11594 5472
rect 11658 5408 11674 5472
rect 11738 5408 11754 5472
rect 11818 5408 11834 5472
rect 11898 5408 11904 5472
rect 12846 5448 13646 5478
rect 11588 5407 11904 5408
rect 841 4994 907 4997
rect 798 4992 907 4994
rect 798 4936 846 4992
rect 902 4936 907 4992
rect 798 4931 907 4936
rect 798 4888 858 4931
rect 0 4798 858 4888
rect 2372 4928 2688 4929
rect 2372 4864 2378 4928
rect 2442 4864 2458 4928
rect 2522 4864 2538 4928
rect 2602 4864 2618 4928
rect 2682 4864 2688 4928
rect 2372 4863 2688 4864
rect 5224 4928 5540 4929
rect 5224 4864 5230 4928
rect 5294 4864 5310 4928
rect 5374 4864 5390 4928
rect 5454 4864 5470 4928
rect 5534 4864 5540 4928
rect 5224 4863 5540 4864
rect 8076 4928 8392 4929
rect 8076 4864 8082 4928
rect 8146 4864 8162 4928
rect 8226 4864 8242 4928
rect 8306 4864 8322 4928
rect 8386 4864 8392 4928
rect 8076 4863 8392 4864
rect 10928 4928 11244 4929
rect 10928 4864 10934 4928
rect 10998 4864 11014 4928
rect 11078 4864 11094 4928
rect 11158 4864 11174 4928
rect 11238 4864 11244 4928
rect 10928 4863 11244 4864
rect 11697 4858 11763 4861
rect 12846 4858 13646 4888
rect 11697 4856 13646 4858
rect 11697 4800 11702 4856
rect 11758 4800 13646 4856
rect 11697 4798 13646 4800
rect 0 4768 800 4798
rect 11697 4795 11763 4798
rect 12846 4768 13646 4798
rect 3032 4384 3348 4385
rect 3032 4320 3038 4384
rect 3102 4320 3118 4384
rect 3182 4320 3198 4384
rect 3262 4320 3278 4384
rect 3342 4320 3348 4384
rect 3032 4319 3348 4320
rect 5884 4384 6200 4385
rect 5884 4320 5890 4384
rect 5954 4320 5970 4384
rect 6034 4320 6050 4384
rect 6114 4320 6130 4384
rect 6194 4320 6200 4384
rect 5884 4319 6200 4320
rect 8736 4384 9052 4385
rect 8736 4320 8742 4384
rect 8806 4320 8822 4384
rect 8886 4320 8902 4384
rect 8966 4320 8982 4384
rect 9046 4320 9052 4384
rect 8736 4319 9052 4320
rect 11588 4384 11904 4385
rect 11588 4320 11594 4384
rect 11658 4320 11674 4384
rect 11738 4320 11754 4384
rect 11818 4320 11834 4384
rect 11898 4320 11904 4384
rect 11588 4319 11904 4320
rect 2372 3840 2688 3841
rect 2372 3776 2378 3840
rect 2442 3776 2458 3840
rect 2522 3776 2538 3840
rect 2602 3776 2618 3840
rect 2682 3776 2688 3840
rect 2372 3775 2688 3776
rect 5224 3840 5540 3841
rect 5224 3776 5230 3840
rect 5294 3776 5310 3840
rect 5374 3776 5390 3840
rect 5454 3776 5470 3840
rect 5534 3776 5540 3840
rect 5224 3775 5540 3776
rect 8076 3840 8392 3841
rect 8076 3776 8082 3840
rect 8146 3776 8162 3840
rect 8226 3776 8242 3840
rect 8306 3776 8322 3840
rect 8386 3776 8392 3840
rect 8076 3775 8392 3776
rect 10928 3840 11244 3841
rect 10928 3776 10934 3840
rect 10998 3776 11014 3840
rect 11078 3776 11094 3840
rect 11158 3776 11174 3840
rect 11238 3776 11244 3840
rect 10928 3775 11244 3776
rect 3032 3296 3348 3297
rect 3032 3232 3038 3296
rect 3102 3232 3118 3296
rect 3182 3232 3198 3296
rect 3262 3232 3278 3296
rect 3342 3232 3348 3296
rect 3032 3231 3348 3232
rect 5884 3296 6200 3297
rect 5884 3232 5890 3296
rect 5954 3232 5970 3296
rect 6034 3232 6050 3296
rect 6114 3232 6130 3296
rect 6194 3232 6200 3296
rect 5884 3231 6200 3232
rect 8736 3296 9052 3297
rect 8736 3232 8742 3296
rect 8806 3232 8822 3296
rect 8886 3232 8902 3296
rect 8966 3232 8982 3296
rect 9046 3232 9052 3296
rect 8736 3231 9052 3232
rect 11588 3296 11904 3297
rect 11588 3232 11594 3296
rect 11658 3232 11674 3296
rect 11738 3232 11754 3296
rect 11818 3232 11834 3296
rect 11898 3232 11904 3296
rect 11588 3231 11904 3232
rect 2372 2752 2688 2753
rect 2372 2688 2378 2752
rect 2442 2688 2458 2752
rect 2522 2688 2538 2752
rect 2602 2688 2618 2752
rect 2682 2688 2688 2752
rect 2372 2687 2688 2688
rect 5224 2752 5540 2753
rect 5224 2688 5230 2752
rect 5294 2688 5310 2752
rect 5374 2688 5390 2752
rect 5454 2688 5470 2752
rect 5534 2688 5540 2752
rect 5224 2687 5540 2688
rect 8076 2752 8392 2753
rect 8076 2688 8082 2752
rect 8146 2688 8162 2752
rect 8226 2688 8242 2752
rect 8306 2688 8322 2752
rect 8386 2688 8392 2752
rect 8076 2687 8392 2688
rect 10928 2752 11244 2753
rect 10928 2688 10934 2752
rect 10998 2688 11014 2752
rect 11078 2688 11094 2752
rect 11158 2688 11174 2752
rect 11238 2688 11244 2752
rect 10928 2687 11244 2688
rect 3032 2208 3348 2209
rect 3032 2144 3038 2208
rect 3102 2144 3118 2208
rect 3182 2144 3198 2208
rect 3262 2144 3278 2208
rect 3342 2144 3348 2208
rect 3032 2143 3348 2144
rect 5884 2208 6200 2209
rect 5884 2144 5890 2208
rect 5954 2144 5970 2208
rect 6034 2144 6050 2208
rect 6114 2144 6130 2208
rect 6194 2144 6200 2208
rect 5884 2143 6200 2144
rect 8736 2208 9052 2209
rect 8736 2144 8742 2208
rect 8806 2144 8822 2208
rect 8886 2144 8902 2208
rect 8966 2144 8982 2208
rect 9046 2144 9052 2208
rect 8736 2143 9052 2144
rect 11588 2208 11904 2209
rect 11588 2144 11594 2208
rect 11658 2144 11674 2208
rect 11738 2144 11754 2208
rect 11818 2144 11834 2208
rect 11898 2144 11904 2208
rect 11588 2143 11904 2144
<< via3 >>
rect 2378 13628 2442 13632
rect 2378 13572 2382 13628
rect 2382 13572 2438 13628
rect 2438 13572 2442 13628
rect 2378 13568 2442 13572
rect 2458 13628 2522 13632
rect 2458 13572 2462 13628
rect 2462 13572 2518 13628
rect 2518 13572 2522 13628
rect 2458 13568 2522 13572
rect 2538 13628 2602 13632
rect 2538 13572 2542 13628
rect 2542 13572 2598 13628
rect 2598 13572 2602 13628
rect 2538 13568 2602 13572
rect 2618 13628 2682 13632
rect 2618 13572 2622 13628
rect 2622 13572 2678 13628
rect 2678 13572 2682 13628
rect 2618 13568 2682 13572
rect 5230 13628 5294 13632
rect 5230 13572 5234 13628
rect 5234 13572 5290 13628
rect 5290 13572 5294 13628
rect 5230 13568 5294 13572
rect 5310 13628 5374 13632
rect 5310 13572 5314 13628
rect 5314 13572 5370 13628
rect 5370 13572 5374 13628
rect 5310 13568 5374 13572
rect 5390 13628 5454 13632
rect 5390 13572 5394 13628
rect 5394 13572 5450 13628
rect 5450 13572 5454 13628
rect 5390 13568 5454 13572
rect 5470 13628 5534 13632
rect 5470 13572 5474 13628
rect 5474 13572 5530 13628
rect 5530 13572 5534 13628
rect 5470 13568 5534 13572
rect 8082 13628 8146 13632
rect 8082 13572 8086 13628
rect 8086 13572 8142 13628
rect 8142 13572 8146 13628
rect 8082 13568 8146 13572
rect 8162 13628 8226 13632
rect 8162 13572 8166 13628
rect 8166 13572 8222 13628
rect 8222 13572 8226 13628
rect 8162 13568 8226 13572
rect 8242 13628 8306 13632
rect 8242 13572 8246 13628
rect 8246 13572 8302 13628
rect 8302 13572 8306 13628
rect 8242 13568 8306 13572
rect 8322 13628 8386 13632
rect 8322 13572 8326 13628
rect 8326 13572 8382 13628
rect 8382 13572 8386 13628
rect 8322 13568 8386 13572
rect 10934 13628 10998 13632
rect 10934 13572 10938 13628
rect 10938 13572 10994 13628
rect 10994 13572 10998 13628
rect 10934 13568 10998 13572
rect 11014 13628 11078 13632
rect 11014 13572 11018 13628
rect 11018 13572 11074 13628
rect 11074 13572 11078 13628
rect 11014 13568 11078 13572
rect 11094 13628 11158 13632
rect 11094 13572 11098 13628
rect 11098 13572 11154 13628
rect 11154 13572 11158 13628
rect 11094 13568 11158 13572
rect 11174 13628 11238 13632
rect 11174 13572 11178 13628
rect 11178 13572 11234 13628
rect 11234 13572 11238 13628
rect 11174 13568 11238 13572
rect 3038 13084 3102 13088
rect 3038 13028 3042 13084
rect 3042 13028 3098 13084
rect 3098 13028 3102 13084
rect 3038 13024 3102 13028
rect 3118 13084 3182 13088
rect 3118 13028 3122 13084
rect 3122 13028 3178 13084
rect 3178 13028 3182 13084
rect 3118 13024 3182 13028
rect 3198 13084 3262 13088
rect 3198 13028 3202 13084
rect 3202 13028 3258 13084
rect 3258 13028 3262 13084
rect 3198 13024 3262 13028
rect 3278 13084 3342 13088
rect 3278 13028 3282 13084
rect 3282 13028 3338 13084
rect 3338 13028 3342 13084
rect 3278 13024 3342 13028
rect 5890 13084 5954 13088
rect 5890 13028 5894 13084
rect 5894 13028 5950 13084
rect 5950 13028 5954 13084
rect 5890 13024 5954 13028
rect 5970 13084 6034 13088
rect 5970 13028 5974 13084
rect 5974 13028 6030 13084
rect 6030 13028 6034 13084
rect 5970 13024 6034 13028
rect 6050 13084 6114 13088
rect 6050 13028 6054 13084
rect 6054 13028 6110 13084
rect 6110 13028 6114 13084
rect 6050 13024 6114 13028
rect 6130 13084 6194 13088
rect 6130 13028 6134 13084
rect 6134 13028 6190 13084
rect 6190 13028 6194 13084
rect 6130 13024 6194 13028
rect 8742 13084 8806 13088
rect 8742 13028 8746 13084
rect 8746 13028 8802 13084
rect 8802 13028 8806 13084
rect 8742 13024 8806 13028
rect 8822 13084 8886 13088
rect 8822 13028 8826 13084
rect 8826 13028 8882 13084
rect 8882 13028 8886 13084
rect 8822 13024 8886 13028
rect 8902 13084 8966 13088
rect 8902 13028 8906 13084
rect 8906 13028 8962 13084
rect 8962 13028 8966 13084
rect 8902 13024 8966 13028
rect 8982 13084 9046 13088
rect 8982 13028 8986 13084
rect 8986 13028 9042 13084
rect 9042 13028 9046 13084
rect 8982 13024 9046 13028
rect 11594 13084 11658 13088
rect 11594 13028 11598 13084
rect 11598 13028 11654 13084
rect 11654 13028 11658 13084
rect 11594 13024 11658 13028
rect 11674 13084 11738 13088
rect 11674 13028 11678 13084
rect 11678 13028 11734 13084
rect 11734 13028 11738 13084
rect 11674 13024 11738 13028
rect 11754 13084 11818 13088
rect 11754 13028 11758 13084
rect 11758 13028 11814 13084
rect 11814 13028 11818 13084
rect 11754 13024 11818 13028
rect 11834 13084 11898 13088
rect 11834 13028 11838 13084
rect 11838 13028 11894 13084
rect 11894 13028 11898 13084
rect 11834 13024 11898 13028
rect 2378 12540 2442 12544
rect 2378 12484 2382 12540
rect 2382 12484 2438 12540
rect 2438 12484 2442 12540
rect 2378 12480 2442 12484
rect 2458 12540 2522 12544
rect 2458 12484 2462 12540
rect 2462 12484 2518 12540
rect 2518 12484 2522 12540
rect 2458 12480 2522 12484
rect 2538 12540 2602 12544
rect 2538 12484 2542 12540
rect 2542 12484 2598 12540
rect 2598 12484 2602 12540
rect 2538 12480 2602 12484
rect 2618 12540 2682 12544
rect 2618 12484 2622 12540
rect 2622 12484 2678 12540
rect 2678 12484 2682 12540
rect 2618 12480 2682 12484
rect 5230 12540 5294 12544
rect 5230 12484 5234 12540
rect 5234 12484 5290 12540
rect 5290 12484 5294 12540
rect 5230 12480 5294 12484
rect 5310 12540 5374 12544
rect 5310 12484 5314 12540
rect 5314 12484 5370 12540
rect 5370 12484 5374 12540
rect 5310 12480 5374 12484
rect 5390 12540 5454 12544
rect 5390 12484 5394 12540
rect 5394 12484 5450 12540
rect 5450 12484 5454 12540
rect 5390 12480 5454 12484
rect 5470 12540 5534 12544
rect 5470 12484 5474 12540
rect 5474 12484 5530 12540
rect 5530 12484 5534 12540
rect 5470 12480 5534 12484
rect 8082 12540 8146 12544
rect 8082 12484 8086 12540
rect 8086 12484 8142 12540
rect 8142 12484 8146 12540
rect 8082 12480 8146 12484
rect 8162 12540 8226 12544
rect 8162 12484 8166 12540
rect 8166 12484 8222 12540
rect 8222 12484 8226 12540
rect 8162 12480 8226 12484
rect 8242 12540 8306 12544
rect 8242 12484 8246 12540
rect 8246 12484 8302 12540
rect 8302 12484 8306 12540
rect 8242 12480 8306 12484
rect 8322 12540 8386 12544
rect 8322 12484 8326 12540
rect 8326 12484 8382 12540
rect 8382 12484 8386 12540
rect 8322 12480 8386 12484
rect 10934 12540 10998 12544
rect 10934 12484 10938 12540
rect 10938 12484 10994 12540
rect 10994 12484 10998 12540
rect 10934 12480 10998 12484
rect 11014 12540 11078 12544
rect 11014 12484 11018 12540
rect 11018 12484 11074 12540
rect 11074 12484 11078 12540
rect 11014 12480 11078 12484
rect 11094 12540 11158 12544
rect 11094 12484 11098 12540
rect 11098 12484 11154 12540
rect 11154 12484 11158 12540
rect 11094 12480 11158 12484
rect 11174 12540 11238 12544
rect 11174 12484 11178 12540
rect 11178 12484 11234 12540
rect 11234 12484 11238 12540
rect 11174 12480 11238 12484
rect 3038 11996 3102 12000
rect 3038 11940 3042 11996
rect 3042 11940 3098 11996
rect 3098 11940 3102 11996
rect 3038 11936 3102 11940
rect 3118 11996 3182 12000
rect 3118 11940 3122 11996
rect 3122 11940 3178 11996
rect 3178 11940 3182 11996
rect 3118 11936 3182 11940
rect 3198 11996 3262 12000
rect 3198 11940 3202 11996
rect 3202 11940 3258 11996
rect 3258 11940 3262 11996
rect 3198 11936 3262 11940
rect 3278 11996 3342 12000
rect 3278 11940 3282 11996
rect 3282 11940 3338 11996
rect 3338 11940 3342 11996
rect 3278 11936 3342 11940
rect 5890 11996 5954 12000
rect 5890 11940 5894 11996
rect 5894 11940 5950 11996
rect 5950 11940 5954 11996
rect 5890 11936 5954 11940
rect 5970 11996 6034 12000
rect 5970 11940 5974 11996
rect 5974 11940 6030 11996
rect 6030 11940 6034 11996
rect 5970 11936 6034 11940
rect 6050 11996 6114 12000
rect 6050 11940 6054 11996
rect 6054 11940 6110 11996
rect 6110 11940 6114 11996
rect 6050 11936 6114 11940
rect 6130 11996 6194 12000
rect 6130 11940 6134 11996
rect 6134 11940 6190 11996
rect 6190 11940 6194 11996
rect 6130 11936 6194 11940
rect 8742 11996 8806 12000
rect 8742 11940 8746 11996
rect 8746 11940 8802 11996
rect 8802 11940 8806 11996
rect 8742 11936 8806 11940
rect 8822 11996 8886 12000
rect 8822 11940 8826 11996
rect 8826 11940 8882 11996
rect 8882 11940 8886 11996
rect 8822 11936 8886 11940
rect 8902 11996 8966 12000
rect 8902 11940 8906 11996
rect 8906 11940 8962 11996
rect 8962 11940 8966 11996
rect 8902 11936 8966 11940
rect 8982 11996 9046 12000
rect 8982 11940 8986 11996
rect 8986 11940 9042 11996
rect 9042 11940 9046 11996
rect 8982 11936 9046 11940
rect 11594 11996 11658 12000
rect 11594 11940 11598 11996
rect 11598 11940 11654 11996
rect 11654 11940 11658 11996
rect 11594 11936 11658 11940
rect 11674 11996 11738 12000
rect 11674 11940 11678 11996
rect 11678 11940 11734 11996
rect 11734 11940 11738 11996
rect 11674 11936 11738 11940
rect 11754 11996 11818 12000
rect 11754 11940 11758 11996
rect 11758 11940 11814 11996
rect 11814 11940 11818 11996
rect 11754 11936 11818 11940
rect 11834 11996 11898 12000
rect 11834 11940 11838 11996
rect 11838 11940 11894 11996
rect 11894 11940 11898 11996
rect 11834 11936 11898 11940
rect 2378 11452 2442 11456
rect 2378 11396 2382 11452
rect 2382 11396 2438 11452
rect 2438 11396 2442 11452
rect 2378 11392 2442 11396
rect 2458 11452 2522 11456
rect 2458 11396 2462 11452
rect 2462 11396 2518 11452
rect 2518 11396 2522 11452
rect 2458 11392 2522 11396
rect 2538 11452 2602 11456
rect 2538 11396 2542 11452
rect 2542 11396 2598 11452
rect 2598 11396 2602 11452
rect 2538 11392 2602 11396
rect 2618 11452 2682 11456
rect 2618 11396 2622 11452
rect 2622 11396 2678 11452
rect 2678 11396 2682 11452
rect 2618 11392 2682 11396
rect 5230 11452 5294 11456
rect 5230 11396 5234 11452
rect 5234 11396 5290 11452
rect 5290 11396 5294 11452
rect 5230 11392 5294 11396
rect 5310 11452 5374 11456
rect 5310 11396 5314 11452
rect 5314 11396 5370 11452
rect 5370 11396 5374 11452
rect 5310 11392 5374 11396
rect 5390 11452 5454 11456
rect 5390 11396 5394 11452
rect 5394 11396 5450 11452
rect 5450 11396 5454 11452
rect 5390 11392 5454 11396
rect 5470 11452 5534 11456
rect 5470 11396 5474 11452
rect 5474 11396 5530 11452
rect 5530 11396 5534 11452
rect 5470 11392 5534 11396
rect 8082 11452 8146 11456
rect 8082 11396 8086 11452
rect 8086 11396 8142 11452
rect 8142 11396 8146 11452
rect 8082 11392 8146 11396
rect 8162 11452 8226 11456
rect 8162 11396 8166 11452
rect 8166 11396 8222 11452
rect 8222 11396 8226 11452
rect 8162 11392 8226 11396
rect 8242 11452 8306 11456
rect 8242 11396 8246 11452
rect 8246 11396 8302 11452
rect 8302 11396 8306 11452
rect 8242 11392 8306 11396
rect 8322 11452 8386 11456
rect 8322 11396 8326 11452
rect 8326 11396 8382 11452
rect 8382 11396 8386 11452
rect 8322 11392 8386 11396
rect 10934 11452 10998 11456
rect 10934 11396 10938 11452
rect 10938 11396 10994 11452
rect 10994 11396 10998 11452
rect 10934 11392 10998 11396
rect 11014 11452 11078 11456
rect 11014 11396 11018 11452
rect 11018 11396 11074 11452
rect 11074 11396 11078 11452
rect 11014 11392 11078 11396
rect 11094 11452 11158 11456
rect 11094 11396 11098 11452
rect 11098 11396 11154 11452
rect 11154 11396 11158 11452
rect 11094 11392 11158 11396
rect 11174 11452 11238 11456
rect 11174 11396 11178 11452
rect 11178 11396 11234 11452
rect 11234 11396 11238 11452
rect 11174 11392 11238 11396
rect 3038 10908 3102 10912
rect 3038 10852 3042 10908
rect 3042 10852 3098 10908
rect 3098 10852 3102 10908
rect 3038 10848 3102 10852
rect 3118 10908 3182 10912
rect 3118 10852 3122 10908
rect 3122 10852 3178 10908
rect 3178 10852 3182 10908
rect 3118 10848 3182 10852
rect 3198 10908 3262 10912
rect 3198 10852 3202 10908
rect 3202 10852 3258 10908
rect 3258 10852 3262 10908
rect 3198 10848 3262 10852
rect 3278 10908 3342 10912
rect 3278 10852 3282 10908
rect 3282 10852 3338 10908
rect 3338 10852 3342 10908
rect 3278 10848 3342 10852
rect 5890 10908 5954 10912
rect 5890 10852 5894 10908
rect 5894 10852 5950 10908
rect 5950 10852 5954 10908
rect 5890 10848 5954 10852
rect 5970 10908 6034 10912
rect 5970 10852 5974 10908
rect 5974 10852 6030 10908
rect 6030 10852 6034 10908
rect 5970 10848 6034 10852
rect 6050 10908 6114 10912
rect 6050 10852 6054 10908
rect 6054 10852 6110 10908
rect 6110 10852 6114 10908
rect 6050 10848 6114 10852
rect 6130 10908 6194 10912
rect 6130 10852 6134 10908
rect 6134 10852 6190 10908
rect 6190 10852 6194 10908
rect 6130 10848 6194 10852
rect 8742 10908 8806 10912
rect 8742 10852 8746 10908
rect 8746 10852 8802 10908
rect 8802 10852 8806 10908
rect 8742 10848 8806 10852
rect 8822 10908 8886 10912
rect 8822 10852 8826 10908
rect 8826 10852 8882 10908
rect 8882 10852 8886 10908
rect 8822 10848 8886 10852
rect 8902 10908 8966 10912
rect 8902 10852 8906 10908
rect 8906 10852 8962 10908
rect 8962 10852 8966 10908
rect 8902 10848 8966 10852
rect 8982 10908 9046 10912
rect 8982 10852 8986 10908
rect 8986 10852 9042 10908
rect 9042 10852 9046 10908
rect 8982 10848 9046 10852
rect 11594 10908 11658 10912
rect 11594 10852 11598 10908
rect 11598 10852 11654 10908
rect 11654 10852 11658 10908
rect 11594 10848 11658 10852
rect 11674 10908 11738 10912
rect 11674 10852 11678 10908
rect 11678 10852 11734 10908
rect 11734 10852 11738 10908
rect 11674 10848 11738 10852
rect 11754 10908 11818 10912
rect 11754 10852 11758 10908
rect 11758 10852 11814 10908
rect 11814 10852 11818 10908
rect 11754 10848 11818 10852
rect 11834 10908 11898 10912
rect 11834 10852 11838 10908
rect 11838 10852 11894 10908
rect 11894 10852 11898 10908
rect 11834 10848 11898 10852
rect 2378 10364 2442 10368
rect 2378 10308 2382 10364
rect 2382 10308 2438 10364
rect 2438 10308 2442 10364
rect 2378 10304 2442 10308
rect 2458 10364 2522 10368
rect 2458 10308 2462 10364
rect 2462 10308 2518 10364
rect 2518 10308 2522 10364
rect 2458 10304 2522 10308
rect 2538 10364 2602 10368
rect 2538 10308 2542 10364
rect 2542 10308 2598 10364
rect 2598 10308 2602 10364
rect 2538 10304 2602 10308
rect 2618 10364 2682 10368
rect 2618 10308 2622 10364
rect 2622 10308 2678 10364
rect 2678 10308 2682 10364
rect 2618 10304 2682 10308
rect 5230 10364 5294 10368
rect 5230 10308 5234 10364
rect 5234 10308 5290 10364
rect 5290 10308 5294 10364
rect 5230 10304 5294 10308
rect 5310 10364 5374 10368
rect 5310 10308 5314 10364
rect 5314 10308 5370 10364
rect 5370 10308 5374 10364
rect 5310 10304 5374 10308
rect 5390 10364 5454 10368
rect 5390 10308 5394 10364
rect 5394 10308 5450 10364
rect 5450 10308 5454 10364
rect 5390 10304 5454 10308
rect 5470 10364 5534 10368
rect 5470 10308 5474 10364
rect 5474 10308 5530 10364
rect 5530 10308 5534 10364
rect 5470 10304 5534 10308
rect 8082 10364 8146 10368
rect 8082 10308 8086 10364
rect 8086 10308 8142 10364
rect 8142 10308 8146 10364
rect 8082 10304 8146 10308
rect 8162 10364 8226 10368
rect 8162 10308 8166 10364
rect 8166 10308 8222 10364
rect 8222 10308 8226 10364
rect 8162 10304 8226 10308
rect 8242 10364 8306 10368
rect 8242 10308 8246 10364
rect 8246 10308 8302 10364
rect 8302 10308 8306 10364
rect 8242 10304 8306 10308
rect 8322 10364 8386 10368
rect 8322 10308 8326 10364
rect 8326 10308 8382 10364
rect 8382 10308 8386 10364
rect 8322 10304 8386 10308
rect 10934 10364 10998 10368
rect 10934 10308 10938 10364
rect 10938 10308 10994 10364
rect 10994 10308 10998 10364
rect 10934 10304 10998 10308
rect 11014 10364 11078 10368
rect 11014 10308 11018 10364
rect 11018 10308 11074 10364
rect 11074 10308 11078 10364
rect 11014 10304 11078 10308
rect 11094 10364 11158 10368
rect 11094 10308 11098 10364
rect 11098 10308 11154 10364
rect 11154 10308 11158 10364
rect 11094 10304 11158 10308
rect 11174 10364 11238 10368
rect 11174 10308 11178 10364
rect 11178 10308 11234 10364
rect 11234 10308 11238 10364
rect 11174 10304 11238 10308
rect 3038 9820 3102 9824
rect 3038 9764 3042 9820
rect 3042 9764 3098 9820
rect 3098 9764 3102 9820
rect 3038 9760 3102 9764
rect 3118 9820 3182 9824
rect 3118 9764 3122 9820
rect 3122 9764 3178 9820
rect 3178 9764 3182 9820
rect 3118 9760 3182 9764
rect 3198 9820 3262 9824
rect 3198 9764 3202 9820
rect 3202 9764 3258 9820
rect 3258 9764 3262 9820
rect 3198 9760 3262 9764
rect 3278 9820 3342 9824
rect 3278 9764 3282 9820
rect 3282 9764 3338 9820
rect 3338 9764 3342 9820
rect 3278 9760 3342 9764
rect 5890 9820 5954 9824
rect 5890 9764 5894 9820
rect 5894 9764 5950 9820
rect 5950 9764 5954 9820
rect 5890 9760 5954 9764
rect 5970 9820 6034 9824
rect 5970 9764 5974 9820
rect 5974 9764 6030 9820
rect 6030 9764 6034 9820
rect 5970 9760 6034 9764
rect 6050 9820 6114 9824
rect 6050 9764 6054 9820
rect 6054 9764 6110 9820
rect 6110 9764 6114 9820
rect 6050 9760 6114 9764
rect 6130 9820 6194 9824
rect 6130 9764 6134 9820
rect 6134 9764 6190 9820
rect 6190 9764 6194 9820
rect 6130 9760 6194 9764
rect 8742 9820 8806 9824
rect 8742 9764 8746 9820
rect 8746 9764 8802 9820
rect 8802 9764 8806 9820
rect 8742 9760 8806 9764
rect 8822 9820 8886 9824
rect 8822 9764 8826 9820
rect 8826 9764 8882 9820
rect 8882 9764 8886 9820
rect 8822 9760 8886 9764
rect 8902 9820 8966 9824
rect 8902 9764 8906 9820
rect 8906 9764 8962 9820
rect 8962 9764 8966 9820
rect 8902 9760 8966 9764
rect 8982 9820 9046 9824
rect 8982 9764 8986 9820
rect 8986 9764 9042 9820
rect 9042 9764 9046 9820
rect 8982 9760 9046 9764
rect 11594 9820 11658 9824
rect 11594 9764 11598 9820
rect 11598 9764 11654 9820
rect 11654 9764 11658 9820
rect 11594 9760 11658 9764
rect 11674 9820 11738 9824
rect 11674 9764 11678 9820
rect 11678 9764 11734 9820
rect 11734 9764 11738 9820
rect 11674 9760 11738 9764
rect 11754 9820 11818 9824
rect 11754 9764 11758 9820
rect 11758 9764 11814 9820
rect 11814 9764 11818 9820
rect 11754 9760 11818 9764
rect 11834 9820 11898 9824
rect 11834 9764 11838 9820
rect 11838 9764 11894 9820
rect 11894 9764 11898 9820
rect 11834 9760 11898 9764
rect 2378 9276 2442 9280
rect 2378 9220 2382 9276
rect 2382 9220 2438 9276
rect 2438 9220 2442 9276
rect 2378 9216 2442 9220
rect 2458 9276 2522 9280
rect 2458 9220 2462 9276
rect 2462 9220 2518 9276
rect 2518 9220 2522 9276
rect 2458 9216 2522 9220
rect 2538 9276 2602 9280
rect 2538 9220 2542 9276
rect 2542 9220 2598 9276
rect 2598 9220 2602 9276
rect 2538 9216 2602 9220
rect 2618 9276 2682 9280
rect 2618 9220 2622 9276
rect 2622 9220 2678 9276
rect 2678 9220 2682 9276
rect 2618 9216 2682 9220
rect 5230 9276 5294 9280
rect 5230 9220 5234 9276
rect 5234 9220 5290 9276
rect 5290 9220 5294 9276
rect 5230 9216 5294 9220
rect 5310 9276 5374 9280
rect 5310 9220 5314 9276
rect 5314 9220 5370 9276
rect 5370 9220 5374 9276
rect 5310 9216 5374 9220
rect 5390 9276 5454 9280
rect 5390 9220 5394 9276
rect 5394 9220 5450 9276
rect 5450 9220 5454 9276
rect 5390 9216 5454 9220
rect 5470 9276 5534 9280
rect 5470 9220 5474 9276
rect 5474 9220 5530 9276
rect 5530 9220 5534 9276
rect 5470 9216 5534 9220
rect 8082 9276 8146 9280
rect 8082 9220 8086 9276
rect 8086 9220 8142 9276
rect 8142 9220 8146 9276
rect 8082 9216 8146 9220
rect 8162 9276 8226 9280
rect 8162 9220 8166 9276
rect 8166 9220 8222 9276
rect 8222 9220 8226 9276
rect 8162 9216 8226 9220
rect 8242 9276 8306 9280
rect 8242 9220 8246 9276
rect 8246 9220 8302 9276
rect 8302 9220 8306 9276
rect 8242 9216 8306 9220
rect 8322 9276 8386 9280
rect 8322 9220 8326 9276
rect 8326 9220 8382 9276
rect 8382 9220 8386 9276
rect 8322 9216 8386 9220
rect 10934 9276 10998 9280
rect 10934 9220 10938 9276
rect 10938 9220 10994 9276
rect 10994 9220 10998 9276
rect 10934 9216 10998 9220
rect 11014 9276 11078 9280
rect 11014 9220 11018 9276
rect 11018 9220 11074 9276
rect 11074 9220 11078 9276
rect 11014 9216 11078 9220
rect 11094 9276 11158 9280
rect 11094 9220 11098 9276
rect 11098 9220 11154 9276
rect 11154 9220 11158 9276
rect 11094 9216 11158 9220
rect 11174 9276 11238 9280
rect 11174 9220 11178 9276
rect 11178 9220 11234 9276
rect 11234 9220 11238 9276
rect 11174 9216 11238 9220
rect 3038 8732 3102 8736
rect 3038 8676 3042 8732
rect 3042 8676 3098 8732
rect 3098 8676 3102 8732
rect 3038 8672 3102 8676
rect 3118 8732 3182 8736
rect 3118 8676 3122 8732
rect 3122 8676 3178 8732
rect 3178 8676 3182 8732
rect 3118 8672 3182 8676
rect 3198 8732 3262 8736
rect 3198 8676 3202 8732
rect 3202 8676 3258 8732
rect 3258 8676 3262 8732
rect 3198 8672 3262 8676
rect 3278 8732 3342 8736
rect 3278 8676 3282 8732
rect 3282 8676 3338 8732
rect 3338 8676 3342 8732
rect 3278 8672 3342 8676
rect 5890 8732 5954 8736
rect 5890 8676 5894 8732
rect 5894 8676 5950 8732
rect 5950 8676 5954 8732
rect 5890 8672 5954 8676
rect 5970 8732 6034 8736
rect 5970 8676 5974 8732
rect 5974 8676 6030 8732
rect 6030 8676 6034 8732
rect 5970 8672 6034 8676
rect 6050 8732 6114 8736
rect 6050 8676 6054 8732
rect 6054 8676 6110 8732
rect 6110 8676 6114 8732
rect 6050 8672 6114 8676
rect 6130 8732 6194 8736
rect 6130 8676 6134 8732
rect 6134 8676 6190 8732
rect 6190 8676 6194 8732
rect 6130 8672 6194 8676
rect 8742 8732 8806 8736
rect 8742 8676 8746 8732
rect 8746 8676 8802 8732
rect 8802 8676 8806 8732
rect 8742 8672 8806 8676
rect 8822 8732 8886 8736
rect 8822 8676 8826 8732
rect 8826 8676 8882 8732
rect 8882 8676 8886 8732
rect 8822 8672 8886 8676
rect 8902 8732 8966 8736
rect 8902 8676 8906 8732
rect 8906 8676 8962 8732
rect 8962 8676 8966 8732
rect 8902 8672 8966 8676
rect 8982 8732 9046 8736
rect 8982 8676 8986 8732
rect 8986 8676 9042 8732
rect 9042 8676 9046 8732
rect 8982 8672 9046 8676
rect 11594 8732 11658 8736
rect 11594 8676 11598 8732
rect 11598 8676 11654 8732
rect 11654 8676 11658 8732
rect 11594 8672 11658 8676
rect 11674 8732 11738 8736
rect 11674 8676 11678 8732
rect 11678 8676 11734 8732
rect 11734 8676 11738 8732
rect 11674 8672 11738 8676
rect 11754 8732 11818 8736
rect 11754 8676 11758 8732
rect 11758 8676 11814 8732
rect 11814 8676 11818 8732
rect 11754 8672 11818 8676
rect 11834 8732 11898 8736
rect 11834 8676 11838 8732
rect 11838 8676 11894 8732
rect 11894 8676 11898 8732
rect 11834 8672 11898 8676
rect 2378 8188 2442 8192
rect 2378 8132 2382 8188
rect 2382 8132 2438 8188
rect 2438 8132 2442 8188
rect 2378 8128 2442 8132
rect 2458 8188 2522 8192
rect 2458 8132 2462 8188
rect 2462 8132 2518 8188
rect 2518 8132 2522 8188
rect 2458 8128 2522 8132
rect 2538 8188 2602 8192
rect 2538 8132 2542 8188
rect 2542 8132 2598 8188
rect 2598 8132 2602 8188
rect 2538 8128 2602 8132
rect 2618 8188 2682 8192
rect 2618 8132 2622 8188
rect 2622 8132 2678 8188
rect 2678 8132 2682 8188
rect 2618 8128 2682 8132
rect 5230 8188 5294 8192
rect 5230 8132 5234 8188
rect 5234 8132 5290 8188
rect 5290 8132 5294 8188
rect 5230 8128 5294 8132
rect 5310 8188 5374 8192
rect 5310 8132 5314 8188
rect 5314 8132 5370 8188
rect 5370 8132 5374 8188
rect 5310 8128 5374 8132
rect 5390 8188 5454 8192
rect 5390 8132 5394 8188
rect 5394 8132 5450 8188
rect 5450 8132 5454 8188
rect 5390 8128 5454 8132
rect 5470 8188 5534 8192
rect 5470 8132 5474 8188
rect 5474 8132 5530 8188
rect 5530 8132 5534 8188
rect 5470 8128 5534 8132
rect 8082 8188 8146 8192
rect 8082 8132 8086 8188
rect 8086 8132 8142 8188
rect 8142 8132 8146 8188
rect 8082 8128 8146 8132
rect 8162 8188 8226 8192
rect 8162 8132 8166 8188
rect 8166 8132 8222 8188
rect 8222 8132 8226 8188
rect 8162 8128 8226 8132
rect 8242 8188 8306 8192
rect 8242 8132 8246 8188
rect 8246 8132 8302 8188
rect 8302 8132 8306 8188
rect 8242 8128 8306 8132
rect 8322 8188 8386 8192
rect 8322 8132 8326 8188
rect 8326 8132 8382 8188
rect 8382 8132 8386 8188
rect 8322 8128 8386 8132
rect 10934 8188 10998 8192
rect 10934 8132 10938 8188
rect 10938 8132 10994 8188
rect 10994 8132 10998 8188
rect 10934 8128 10998 8132
rect 11014 8188 11078 8192
rect 11014 8132 11018 8188
rect 11018 8132 11074 8188
rect 11074 8132 11078 8188
rect 11014 8128 11078 8132
rect 11094 8188 11158 8192
rect 11094 8132 11098 8188
rect 11098 8132 11154 8188
rect 11154 8132 11158 8188
rect 11094 8128 11158 8132
rect 11174 8188 11238 8192
rect 11174 8132 11178 8188
rect 11178 8132 11234 8188
rect 11234 8132 11238 8188
rect 11174 8128 11238 8132
rect 3038 7644 3102 7648
rect 3038 7588 3042 7644
rect 3042 7588 3098 7644
rect 3098 7588 3102 7644
rect 3038 7584 3102 7588
rect 3118 7644 3182 7648
rect 3118 7588 3122 7644
rect 3122 7588 3178 7644
rect 3178 7588 3182 7644
rect 3118 7584 3182 7588
rect 3198 7644 3262 7648
rect 3198 7588 3202 7644
rect 3202 7588 3258 7644
rect 3258 7588 3262 7644
rect 3198 7584 3262 7588
rect 3278 7644 3342 7648
rect 3278 7588 3282 7644
rect 3282 7588 3338 7644
rect 3338 7588 3342 7644
rect 3278 7584 3342 7588
rect 5890 7644 5954 7648
rect 5890 7588 5894 7644
rect 5894 7588 5950 7644
rect 5950 7588 5954 7644
rect 5890 7584 5954 7588
rect 5970 7644 6034 7648
rect 5970 7588 5974 7644
rect 5974 7588 6030 7644
rect 6030 7588 6034 7644
rect 5970 7584 6034 7588
rect 6050 7644 6114 7648
rect 6050 7588 6054 7644
rect 6054 7588 6110 7644
rect 6110 7588 6114 7644
rect 6050 7584 6114 7588
rect 6130 7644 6194 7648
rect 6130 7588 6134 7644
rect 6134 7588 6190 7644
rect 6190 7588 6194 7644
rect 6130 7584 6194 7588
rect 8742 7644 8806 7648
rect 8742 7588 8746 7644
rect 8746 7588 8802 7644
rect 8802 7588 8806 7644
rect 8742 7584 8806 7588
rect 8822 7644 8886 7648
rect 8822 7588 8826 7644
rect 8826 7588 8882 7644
rect 8882 7588 8886 7644
rect 8822 7584 8886 7588
rect 8902 7644 8966 7648
rect 8902 7588 8906 7644
rect 8906 7588 8962 7644
rect 8962 7588 8966 7644
rect 8902 7584 8966 7588
rect 8982 7644 9046 7648
rect 8982 7588 8986 7644
rect 8986 7588 9042 7644
rect 9042 7588 9046 7644
rect 8982 7584 9046 7588
rect 11594 7644 11658 7648
rect 11594 7588 11598 7644
rect 11598 7588 11654 7644
rect 11654 7588 11658 7644
rect 11594 7584 11658 7588
rect 11674 7644 11738 7648
rect 11674 7588 11678 7644
rect 11678 7588 11734 7644
rect 11734 7588 11738 7644
rect 11674 7584 11738 7588
rect 11754 7644 11818 7648
rect 11754 7588 11758 7644
rect 11758 7588 11814 7644
rect 11814 7588 11818 7644
rect 11754 7584 11818 7588
rect 11834 7644 11898 7648
rect 11834 7588 11838 7644
rect 11838 7588 11894 7644
rect 11894 7588 11898 7644
rect 11834 7584 11898 7588
rect 2378 7100 2442 7104
rect 2378 7044 2382 7100
rect 2382 7044 2438 7100
rect 2438 7044 2442 7100
rect 2378 7040 2442 7044
rect 2458 7100 2522 7104
rect 2458 7044 2462 7100
rect 2462 7044 2518 7100
rect 2518 7044 2522 7100
rect 2458 7040 2522 7044
rect 2538 7100 2602 7104
rect 2538 7044 2542 7100
rect 2542 7044 2598 7100
rect 2598 7044 2602 7100
rect 2538 7040 2602 7044
rect 2618 7100 2682 7104
rect 2618 7044 2622 7100
rect 2622 7044 2678 7100
rect 2678 7044 2682 7100
rect 2618 7040 2682 7044
rect 5230 7100 5294 7104
rect 5230 7044 5234 7100
rect 5234 7044 5290 7100
rect 5290 7044 5294 7100
rect 5230 7040 5294 7044
rect 5310 7100 5374 7104
rect 5310 7044 5314 7100
rect 5314 7044 5370 7100
rect 5370 7044 5374 7100
rect 5310 7040 5374 7044
rect 5390 7100 5454 7104
rect 5390 7044 5394 7100
rect 5394 7044 5450 7100
rect 5450 7044 5454 7100
rect 5390 7040 5454 7044
rect 5470 7100 5534 7104
rect 5470 7044 5474 7100
rect 5474 7044 5530 7100
rect 5530 7044 5534 7100
rect 5470 7040 5534 7044
rect 8082 7100 8146 7104
rect 8082 7044 8086 7100
rect 8086 7044 8142 7100
rect 8142 7044 8146 7100
rect 8082 7040 8146 7044
rect 8162 7100 8226 7104
rect 8162 7044 8166 7100
rect 8166 7044 8222 7100
rect 8222 7044 8226 7100
rect 8162 7040 8226 7044
rect 8242 7100 8306 7104
rect 8242 7044 8246 7100
rect 8246 7044 8302 7100
rect 8302 7044 8306 7100
rect 8242 7040 8306 7044
rect 8322 7100 8386 7104
rect 8322 7044 8326 7100
rect 8326 7044 8382 7100
rect 8382 7044 8386 7100
rect 8322 7040 8386 7044
rect 10934 7100 10998 7104
rect 10934 7044 10938 7100
rect 10938 7044 10994 7100
rect 10994 7044 10998 7100
rect 10934 7040 10998 7044
rect 11014 7100 11078 7104
rect 11014 7044 11018 7100
rect 11018 7044 11074 7100
rect 11074 7044 11078 7100
rect 11014 7040 11078 7044
rect 11094 7100 11158 7104
rect 11094 7044 11098 7100
rect 11098 7044 11154 7100
rect 11154 7044 11158 7100
rect 11094 7040 11158 7044
rect 11174 7100 11238 7104
rect 11174 7044 11178 7100
rect 11178 7044 11234 7100
rect 11234 7044 11238 7100
rect 11174 7040 11238 7044
rect 3038 6556 3102 6560
rect 3038 6500 3042 6556
rect 3042 6500 3098 6556
rect 3098 6500 3102 6556
rect 3038 6496 3102 6500
rect 3118 6556 3182 6560
rect 3118 6500 3122 6556
rect 3122 6500 3178 6556
rect 3178 6500 3182 6556
rect 3118 6496 3182 6500
rect 3198 6556 3262 6560
rect 3198 6500 3202 6556
rect 3202 6500 3258 6556
rect 3258 6500 3262 6556
rect 3198 6496 3262 6500
rect 3278 6556 3342 6560
rect 3278 6500 3282 6556
rect 3282 6500 3338 6556
rect 3338 6500 3342 6556
rect 3278 6496 3342 6500
rect 5890 6556 5954 6560
rect 5890 6500 5894 6556
rect 5894 6500 5950 6556
rect 5950 6500 5954 6556
rect 5890 6496 5954 6500
rect 5970 6556 6034 6560
rect 5970 6500 5974 6556
rect 5974 6500 6030 6556
rect 6030 6500 6034 6556
rect 5970 6496 6034 6500
rect 6050 6556 6114 6560
rect 6050 6500 6054 6556
rect 6054 6500 6110 6556
rect 6110 6500 6114 6556
rect 6050 6496 6114 6500
rect 6130 6556 6194 6560
rect 6130 6500 6134 6556
rect 6134 6500 6190 6556
rect 6190 6500 6194 6556
rect 6130 6496 6194 6500
rect 8742 6556 8806 6560
rect 8742 6500 8746 6556
rect 8746 6500 8802 6556
rect 8802 6500 8806 6556
rect 8742 6496 8806 6500
rect 8822 6556 8886 6560
rect 8822 6500 8826 6556
rect 8826 6500 8882 6556
rect 8882 6500 8886 6556
rect 8822 6496 8886 6500
rect 8902 6556 8966 6560
rect 8902 6500 8906 6556
rect 8906 6500 8962 6556
rect 8962 6500 8966 6556
rect 8902 6496 8966 6500
rect 8982 6556 9046 6560
rect 8982 6500 8986 6556
rect 8986 6500 9042 6556
rect 9042 6500 9046 6556
rect 8982 6496 9046 6500
rect 11594 6556 11658 6560
rect 11594 6500 11598 6556
rect 11598 6500 11654 6556
rect 11654 6500 11658 6556
rect 11594 6496 11658 6500
rect 11674 6556 11738 6560
rect 11674 6500 11678 6556
rect 11678 6500 11734 6556
rect 11734 6500 11738 6556
rect 11674 6496 11738 6500
rect 11754 6556 11818 6560
rect 11754 6500 11758 6556
rect 11758 6500 11814 6556
rect 11814 6500 11818 6556
rect 11754 6496 11818 6500
rect 11834 6556 11898 6560
rect 11834 6500 11838 6556
rect 11838 6500 11894 6556
rect 11894 6500 11898 6556
rect 11834 6496 11898 6500
rect 2378 6012 2442 6016
rect 2378 5956 2382 6012
rect 2382 5956 2438 6012
rect 2438 5956 2442 6012
rect 2378 5952 2442 5956
rect 2458 6012 2522 6016
rect 2458 5956 2462 6012
rect 2462 5956 2518 6012
rect 2518 5956 2522 6012
rect 2458 5952 2522 5956
rect 2538 6012 2602 6016
rect 2538 5956 2542 6012
rect 2542 5956 2598 6012
rect 2598 5956 2602 6012
rect 2538 5952 2602 5956
rect 2618 6012 2682 6016
rect 2618 5956 2622 6012
rect 2622 5956 2678 6012
rect 2678 5956 2682 6012
rect 2618 5952 2682 5956
rect 5230 6012 5294 6016
rect 5230 5956 5234 6012
rect 5234 5956 5290 6012
rect 5290 5956 5294 6012
rect 5230 5952 5294 5956
rect 5310 6012 5374 6016
rect 5310 5956 5314 6012
rect 5314 5956 5370 6012
rect 5370 5956 5374 6012
rect 5310 5952 5374 5956
rect 5390 6012 5454 6016
rect 5390 5956 5394 6012
rect 5394 5956 5450 6012
rect 5450 5956 5454 6012
rect 5390 5952 5454 5956
rect 5470 6012 5534 6016
rect 5470 5956 5474 6012
rect 5474 5956 5530 6012
rect 5530 5956 5534 6012
rect 5470 5952 5534 5956
rect 8082 6012 8146 6016
rect 8082 5956 8086 6012
rect 8086 5956 8142 6012
rect 8142 5956 8146 6012
rect 8082 5952 8146 5956
rect 8162 6012 8226 6016
rect 8162 5956 8166 6012
rect 8166 5956 8222 6012
rect 8222 5956 8226 6012
rect 8162 5952 8226 5956
rect 8242 6012 8306 6016
rect 8242 5956 8246 6012
rect 8246 5956 8302 6012
rect 8302 5956 8306 6012
rect 8242 5952 8306 5956
rect 8322 6012 8386 6016
rect 8322 5956 8326 6012
rect 8326 5956 8382 6012
rect 8382 5956 8386 6012
rect 8322 5952 8386 5956
rect 10934 6012 10998 6016
rect 10934 5956 10938 6012
rect 10938 5956 10994 6012
rect 10994 5956 10998 6012
rect 10934 5952 10998 5956
rect 11014 6012 11078 6016
rect 11014 5956 11018 6012
rect 11018 5956 11074 6012
rect 11074 5956 11078 6012
rect 11014 5952 11078 5956
rect 11094 6012 11158 6016
rect 11094 5956 11098 6012
rect 11098 5956 11154 6012
rect 11154 5956 11158 6012
rect 11094 5952 11158 5956
rect 11174 6012 11238 6016
rect 11174 5956 11178 6012
rect 11178 5956 11234 6012
rect 11234 5956 11238 6012
rect 11174 5952 11238 5956
rect 3038 5468 3102 5472
rect 3038 5412 3042 5468
rect 3042 5412 3098 5468
rect 3098 5412 3102 5468
rect 3038 5408 3102 5412
rect 3118 5468 3182 5472
rect 3118 5412 3122 5468
rect 3122 5412 3178 5468
rect 3178 5412 3182 5468
rect 3118 5408 3182 5412
rect 3198 5468 3262 5472
rect 3198 5412 3202 5468
rect 3202 5412 3258 5468
rect 3258 5412 3262 5468
rect 3198 5408 3262 5412
rect 3278 5468 3342 5472
rect 3278 5412 3282 5468
rect 3282 5412 3338 5468
rect 3338 5412 3342 5468
rect 3278 5408 3342 5412
rect 5890 5468 5954 5472
rect 5890 5412 5894 5468
rect 5894 5412 5950 5468
rect 5950 5412 5954 5468
rect 5890 5408 5954 5412
rect 5970 5468 6034 5472
rect 5970 5412 5974 5468
rect 5974 5412 6030 5468
rect 6030 5412 6034 5468
rect 5970 5408 6034 5412
rect 6050 5468 6114 5472
rect 6050 5412 6054 5468
rect 6054 5412 6110 5468
rect 6110 5412 6114 5468
rect 6050 5408 6114 5412
rect 6130 5468 6194 5472
rect 6130 5412 6134 5468
rect 6134 5412 6190 5468
rect 6190 5412 6194 5468
rect 6130 5408 6194 5412
rect 8742 5468 8806 5472
rect 8742 5412 8746 5468
rect 8746 5412 8802 5468
rect 8802 5412 8806 5468
rect 8742 5408 8806 5412
rect 8822 5468 8886 5472
rect 8822 5412 8826 5468
rect 8826 5412 8882 5468
rect 8882 5412 8886 5468
rect 8822 5408 8886 5412
rect 8902 5468 8966 5472
rect 8902 5412 8906 5468
rect 8906 5412 8962 5468
rect 8962 5412 8966 5468
rect 8902 5408 8966 5412
rect 8982 5468 9046 5472
rect 8982 5412 8986 5468
rect 8986 5412 9042 5468
rect 9042 5412 9046 5468
rect 8982 5408 9046 5412
rect 11594 5468 11658 5472
rect 11594 5412 11598 5468
rect 11598 5412 11654 5468
rect 11654 5412 11658 5468
rect 11594 5408 11658 5412
rect 11674 5468 11738 5472
rect 11674 5412 11678 5468
rect 11678 5412 11734 5468
rect 11734 5412 11738 5468
rect 11674 5408 11738 5412
rect 11754 5468 11818 5472
rect 11754 5412 11758 5468
rect 11758 5412 11814 5468
rect 11814 5412 11818 5468
rect 11754 5408 11818 5412
rect 11834 5468 11898 5472
rect 11834 5412 11838 5468
rect 11838 5412 11894 5468
rect 11894 5412 11898 5468
rect 11834 5408 11898 5412
rect 2378 4924 2442 4928
rect 2378 4868 2382 4924
rect 2382 4868 2438 4924
rect 2438 4868 2442 4924
rect 2378 4864 2442 4868
rect 2458 4924 2522 4928
rect 2458 4868 2462 4924
rect 2462 4868 2518 4924
rect 2518 4868 2522 4924
rect 2458 4864 2522 4868
rect 2538 4924 2602 4928
rect 2538 4868 2542 4924
rect 2542 4868 2598 4924
rect 2598 4868 2602 4924
rect 2538 4864 2602 4868
rect 2618 4924 2682 4928
rect 2618 4868 2622 4924
rect 2622 4868 2678 4924
rect 2678 4868 2682 4924
rect 2618 4864 2682 4868
rect 5230 4924 5294 4928
rect 5230 4868 5234 4924
rect 5234 4868 5290 4924
rect 5290 4868 5294 4924
rect 5230 4864 5294 4868
rect 5310 4924 5374 4928
rect 5310 4868 5314 4924
rect 5314 4868 5370 4924
rect 5370 4868 5374 4924
rect 5310 4864 5374 4868
rect 5390 4924 5454 4928
rect 5390 4868 5394 4924
rect 5394 4868 5450 4924
rect 5450 4868 5454 4924
rect 5390 4864 5454 4868
rect 5470 4924 5534 4928
rect 5470 4868 5474 4924
rect 5474 4868 5530 4924
rect 5530 4868 5534 4924
rect 5470 4864 5534 4868
rect 8082 4924 8146 4928
rect 8082 4868 8086 4924
rect 8086 4868 8142 4924
rect 8142 4868 8146 4924
rect 8082 4864 8146 4868
rect 8162 4924 8226 4928
rect 8162 4868 8166 4924
rect 8166 4868 8222 4924
rect 8222 4868 8226 4924
rect 8162 4864 8226 4868
rect 8242 4924 8306 4928
rect 8242 4868 8246 4924
rect 8246 4868 8302 4924
rect 8302 4868 8306 4924
rect 8242 4864 8306 4868
rect 8322 4924 8386 4928
rect 8322 4868 8326 4924
rect 8326 4868 8382 4924
rect 8382 4868 8386 4924
rect 8322 4864 8386 4868
rect 10934 4924 10998 4928
rect 10934 4868 10938 4924
rect 10938 4868 10994 4924
rect 10994 4868 10998 4924
rect 10934 4864 10998 4868
rect 11014 4924 11078 4928
rect 11014 4868 11018 4924
rect 11018 4868 11074 4924
rect 11074 4868 11078 4924
rect 11014 4864 11078 4868
rect 11094 4924 11158 4928
rect 11094 4868 11098 4924
rect 11098 4868 11154 4924
rect 11154 4868 11158 4924
rect 11094 4864 11158 4868
rect 11174 4924 11238 4928
rect 11174 4868 11178 4924
rect 11178 4868 11234 4924
rect 11234 4868 11238 4924
rect 11174 4864 11238 4868
rect 3038 4380 3102 4384
rect 3038 4324 3042 4380
rect 3042 4324 3098 4380
rect 3098 4324 3102 4380
rect 3038 4320 3102 4324
rect 3118 4380 3182 4384
rect 3118 4324 3122 4380
rect 3122 4324 3178 4380
rect 3178 4324 3182 4380
rect 3118 4320 3182 4324
rect 3198 4380 3262 4384
rect 3198 4324 3202 4380
rect 3202 4324 3258 4380
rect 3258 4324 3262 4380
rect 3198 4320 3262 4324
rect 3278 4380 3342 4384
rect 3278 4324 3282 4380
rect 3282 4324 3338 4380
rect 3338 4324 3342 4380
rect 3278 4320 3342 4324
rect 5890 4380 5954 4384
rect 5890 4324 5894 4380
rect 5894 4324 5950 4380
rect 5950 4324 5954 4380
rect 5890 4320 5954 4324
rect 5970 4380 6034 4384
rect 5970 4324 5974 4380
rect 5974 4324 6030 4380
rect 6030 4324 6034 4380
rect 5970 4320 6034 4324
rect 6050 4380 6114 4384
rect 6050 4324 6054 4380
rect 6054 4324 6110 4380
rect 6110 4324 6114 4380
rect 6050 4320 6114 4324
rect 6130 4380 6194 4384
rect 6130 4324 6134 4380
rect 6134 4324 6190 4380
rect 6190 4324 6194 4380
rect 6130 4320 6194 4324
rect 8742 4380 8806 4384
rect 8742 4324 8746 4380
rect 8746 4324 8802 4380
rect 8802 4324 8806 4380
rect 8742 4320 8806 4324
rect 8822 4380 8886 4384
rect 8822 4324 8826 4380
rect 8826 4324 8882 4380
rect 8882 4324 8886 4380
rect 8822 4320 8886 4324
rect 8902 4380 8966 4384
rect 8902 4324 8906 4380
rect 8906 4324 8962 4380
rect 8962 4324 8966 4380
rect 8902 4320 8966 4324
rect 8982 4380 9046 4384
rect 8982 4324 8986 4380
rect 8986 4324 9042 4380
rect 9042 4324 9046 4380
rect 8982 4320 9046 4324
rect 11594 4380 11658 4384
rect 11594 4324 11598 4380
rect 11598 4324 11654 4380
rect 11654 4324 11658 4380
rect 11594 4320 11658 4324
rect 11674 4380 11738 4384
rect 11674 4324 11678 4380
rect 11678 4324 11734 4380
rect 11734 4324 11738 4380
rect 11674 4320 11738 4324
rect 11754 4380 11818 4384
rect 11754 4324 11758 4380
rect 11758 4324 11814 4380
rect 11814 4324 11818 4380
rect 11754 4320 11818 4324
rect 11834 4380 11898 4384
rect 11834 4324 11838 4380
rect 11838 4324 11894 4380
rect 11894 4324 11898 4380
rect 11834 4320 11898 4324
rect 2378 3836 2442 3840
rect 2378 3780 2382 3836
rect 2382 3780 2438 3836
rect 2438 3780 2442 3836
rect 2378 3776 2442 3780
rect 2458 3836 2522 3840
rect 2458 3780 2462 3836
rect 2462 3780 2518 3836
rect 2518 3780 2522 3836
rect 2458 3776 2522 3780
rect 2538 3836 2602 3840
rect 2538 3780 2542 3836
rect 2542 3780 2598 3836
rect 2598 3780 2602 3836
rect 2538 3776 2602 3780
rect 2618 3836 2682 3840
rect 2618 3780 2622 3836
rect 2622 3780 2678 3836
rect 2678 3780 2682 3836
rect 2618 3776 2682 3780
rect 5230 3836 5294 3840
rect 5230 3780 5234 3836
rect 5234 3780 5290 3836
rect 5290 3780 5294 3836
rect 5230 3776 5294 3780
rect 5310 3836 5374 3840
rect 5310 3780 5314 3836
rect 5314 3780 5370 3836
rect 5370 3780 5374 3836
rect 5310 3776 5374 3780
rect 5390 3836 5454 3840
rect 5390 3780 5394 3836
rect 5394 3780 5450 3836
rect 5450 3780 5454 3836
rect 5390 3776 5454 3780
rect 5470 3836 5534 3840
rect 5470 3780 5474 3836
rect 5474 3780 5530 3836
rect 5530 3780 5534 3836
rect 5470 3776 5534 3780
rect 8082 3836 8146 3840
rect 8082 3780 8086 3836
rect 8086 3780 8142 3836
rect 8142 3780 8146 3836
rect 8082 3776 8146 3780
rect 8162 3836 8226 3840
rect 8162 3780 8166 3836
rect 8166 3780 8222 3836
rect 8222 3780 8226 3836
rect 8162 3776 8226 3780
rect 8242 3836 8306 3840
rect 8242 3780 8246 3836
rect 8246 3780 8302 3836
rect 8302 3780 8306 3836
rect 8242 3776 8306 3780
rect 8322 3836 8386 3840
rect 8322 3780 8326 3836
rect 8326 3780 8382 3836
rect 8382 3780 8386 3836
rect 8322 3776 8386 3780
rect 10934 3836 10998 3840
rect 10934 3780 10938 3836
rect 10938 3780 10994 3836
rect 10994 3780 10998 3836
rect 10934 3776 10998 3780
rect 11014 3836 11078 3840
rect 11014 3780 11018 3836
rect 11018 3780 11074 3836
rect 11074 3780 11078 3836
rect 11014 3776 11078 3780
rect 11094 3836 11158 3840
rect 11094 3780 11098 3836
rect 11098 3780 11154 3836
rect 11154 3780 11158 3836
rect 11094 3776 11158 3780
rect 11174 3836 11238 3840
rect 11174 3780 11178 3836
rect 11178 3780 11234 3836
rect 11234 3780 11238 3836
rect 11174 3776 11238 3780
rect 3038 3292 3102 3296
rect 3038 3236 3042 3292
rect 3042 3236 3098 3292
rect 3098 3236 3102 3292
rect 3038 3232 3102 3236
rect 3118 3292 3182 3296
rect 3118 3236 3122 3292
rect 3122 3236 3178 3292
rect 3178 3236 3182 3292
rect 3118 3232 3182 3236
rect 3198 3292 3262 3296
rect 3198 3236 3202 3292
rect 3202 3236 3258 3292
rect 3258 3236 3262 3292
rect 3198 3232 3262 3236
rect 3278 3292 3342 3296
rect 3278 3236 3282 3292
rect 3282 3236 3338 3292
rect 3338 3236 3342 3292
rect 3278 3232 3342 3236
rect 5890 3292 5954 3296
rect 5890 3236 5894 3292
rect 5894 3236 5950 3292
rect 5950 3236 5954 3292
rect 5890 3232 5954 3236
rect 5970 3292 6034 3296
rect 5970 3236 5974 3292
rect 5974 3236 6030 3292
rect 6030 3236 6034 3292
rect 5970 3232 6034 3236
rect 6050 3292 6114 3296
rect 6050 3236 6054 3292
rect 6054 3236 6110 3292
rect 6110 3236 6114 3292
rect 6050 3232 6114 3236
rect 6130 3292 6194 3296
rect 6130 3236 6134 3292
rect 6134 3236 6190 3292
rect 6190 3236 6194 3292
rect 6130 3232 6194 3236
rect 8742 3292 8806 3296
rect 8742 3236 8746 3292
rect 8746 3236 8802 3292
rect 8802 3236 8806 3292
rect 8742 3232 8806 3236
rect 8822 3292 8886 3296
rect 8822 3236 8826 3292
rect 8826 3236 8882 3292
rect 8882 3236 8886 3292
rect 8822 3232 8886 3236
rect 8902 3292 8966 3296
rect 8902 3236 8906 3292
rect 8906 3236 8962 3292
rect 8962 3236 8966 3292
rect 8902 3232 8966 3236
rect 8982 3292 9046 3296
rect 8982 3236 8986 3292
rect 8986 3236 9042 3292
rect 9042 3236 9046 3292
rect 8982 3232 9046 3236
rect 11594 3292 11658 3296
rect 11594 3236 11598 3292
rect 11598 3236 11654 3292
rect 11654 3236 11658 3292
rect 11594 3232 11658 3236
rect 11674 3292 11738 3296
rect 11674 3236 11678 3292
rect 11678 3236 11734 3292
rect 11734 3236 11738 3292
rect 11674 3232 11738 3236
rect 11754 3292 11818 3296
rect 11754 3236 11758 3292
rect 11758 3236 11814 3292
rect 11814 3236 11818 3292
rect 11754 3232 11818 3236
rect 11834 3292 11898 3296
rect 11834 3236 11838 3292
rect 11838 3236 11894 3292
rect 11894 3236 11898 3292
rect 11834 3232 11898 3236
rect 2378 2748 2442 2752
rect 2378 2692 2382 2748
rect 2382 2692 2438 2748
rect 2438 2692 2442 2748
rect 2378 2688 2442 2692
rect 2458 2748 2522 2752
rect 2458 2692 2462 2748
rect 2462 2692 2518 2748
rect 2518 2692 2522 2748
rect 2458 2688 2522 2692
rect 2538 2748 2602 2752
rect 2538 2692 2542 2748
rect 2542 2692 2598 2748
rect 2598 2692 2602 2748
rect 2538 2688 2602 2692
rect 2618 2748 2682 2752
rect 2618 2692 2622 2748
rect 2622 2692 2678 2748
rect 2678 2692 2682 2748
rect 2618 2688 2682 2692
rect 5230 2748 5294 2752
rect 5230 2692 5234 2748
rect 5234 2692 5290 2748
rect 5290 2692 5294 2748
rect 5230 2688 5294 2692
rect 5310 2748 5374 2752
rect 5310 2692 5314 2748
rect 5314 2692 5370 2748
rect 5370 2692 5374 2748
rect 5310 2688 5374 2692
rect 5390 2748 5454 2752
rect 5390 2692 5394 2748
rect 5394 2692 5450 2748
rect 5450 2692 5454 2748
rect 5390 2688 5454 2692
rect 5470 2748 5534 2752
rect 5470 2692 5474 2748
rect 5474 2692 5530 2748
rect 5530 2692 5534 2748
rect 5470 2688 5534 2692
rect 8082 2748 8146 2752
rect 8082 2692 8086 2748
rect 8086 2692 8142 2748
rect 8142 2692 8146 2748
rect 8082 2688 8146 2692
rect 8162 2748 8226 2752
rect 8162 2692 8166 2748
rect 8166 2692 8222 2748
rect 8222 2692 8226 2748
rect 8162 2688 8226 2692
rect 8242 2748 8306 2752
rect 8242 2692 8246 2748
rect 8246 2692 8302 2748
rect 8302 2692 8306 2748
rect 8242 2688 8306 2692
rect 8322 2748 8386 2752
rect 8322 2692 8326 2748
rect 8326 2692 8382 2748
rect 8382 2692 8386 2748
rect 8322 2688 8386 2692
rect 10934 2748 10998 2752
rect 10934 2692 10938 2748
rect 10938 2692 10994 2748
rect 10994 2692 10998 2748
rect 10934 2688 10998 2692
rect 11014 2748 11078 2752
rect 11014 2692 11018 2748
rect 11018 2692 11074 2748
rect 11074 2692 11078 2748
rect 11014 2688 11078 2692
rect 11094 2748 11158 2752
rect 11094 2692 11098 2748
rect 11098 2692 11154 2748
rect 11154 2692 11158 2748
rect 11094 2688 11158 2692
rect 11174 2748 11238 2752
rect 11174 2692 11178 2748
rect 11178 2692 11234 2748
rect 11234 2692 11238 2748
rect 11174 2688 11238 2692
rect 3038 2204 3102 2208
rect 3038 2148 3042 2204
rect 3042 2148 3098 2204
rect 3098 2148 3102 2204
rect 3038 2144 3102 2148
rect 3118 2204 3182 2208
rect 3118 2148 3122 2204
rect 3122 2148 3178 2204
rect 3178 2148 3182 2204
rect 3118 2144 3182 2148
rect 3198 2204 3262 2208
rect 3198 2148 3202 2204
rect 3202 2148 3258 2204
rect 3258 2148 3262 2204
rect 3198 2144 3262 2148
rect 3278 2204 3342 2208
rect 3278 2148 3282 2204
rect 3282 2148 3338 2204
rect 3338 2148 3342 2204
rect 3278 2144 3342 2148
rect 5890 2204 5954 2208
rect 5890 2148 5894 2204
rect 5894 2148 5950 2204
rect 5950 2148 5954 2204
rect 5890 2144 5954 2148
rect 5970 2204 6034 2208
rect 5970 2148 5974 2204
rect 5974 2148 6030 2204
rect 6030 2148 6034 2204
rect 5970 2144 6034 2148
rect 6050 2204 6114 2208
rect 6050 2148 6054 2204
rect 6054 2148 6110 2204
rect 6110 2148 6114 2204
rect 6050 2144 6114 2148
rect 6130 2204 6194 2208
rect 6130 2148 6134 2204
rect 6134 2148 6190 2204
rect 6190 2148 6194 2204
rect 6130 2144 6194 2148
rect 8742 2204 8806 2208
rect 8742 2148 8746 2204
rect 8746 2148 8802 2204
rect 8802 2148 8806 2204
rect 8742 2144 8806 2148
rect 8822 2204 8886 2208
rect 8822 2148 8826 2204
rect 8826 2148 8882 2204
rect 8882 2148 8886 2204
rect 8822 2144 8886 2148
rect 8902 2204 8966 2208
rect 8902 2148 8906 2204
rect 8906 2148 8962 2204
rect 8962 2148 8966 2204
rect 8902 2144 8966 2148
rect 8982 2204 9046 2208
rect 8982 2148 8986 2204
rect 8986 2148 9042 2204
rect 9042 2148 9046 2204
rect 8982 2144 9046 2148
rect 11594 2204 11658 2208
rect 11594 2148 11598 2204
rect 11598 2148 11654 2204
rect 11654 2148 11658 2204
rect 11594 2144 11658 2148
rect 11674 2204 11738 2208
rect 11674 2148 11678 2204
rect 11678 2148 11734 2204
rect 11734 2148 11738 2204
rect 11674 2144 11738 2148
rect 11754 2204 11818 2208
rect 11754 2148 11758 2204
rect 11758 2148 11814 2204
rect 11814 2148 11818 2204
rect 11754 2144 11818 2148
rect 11834 2204 11898 2208
rect 11834 2148 11838 2204
rect 11838 2148 11894 2204
rect 11894 2148 11898 2204
rect 11834 2144 11898 2148
<< metal4 >>
rect 2370 13632 2690 13648
rect 2370 13568 2378 13632
rect 2442 13568 2458 13632
rect 2522 13568 2538 13632
rect 2602 13568 2618 13632
rect 2682 13568 2690 13632
rect 2370 12544 2690 13568
rect 2370 12480 2378 12544
rect 2442 12480 2458 12544
rect 2522 12480 2538 12544
rect 2602 12480 2618 12544
rect 2682 12480 2690 12544
rect 2370 12290 2690 12480
rect 2370 12054 2412 12290
rect 2648 12054 2690 12290
rect 2370 11456 2690 12054
rect 2370 11392 2378 11456
rect 2442 11392 2458 11456
rect 2522 11392 2538 11456
rect 2602 11392 2618 11456
rect 2682 11392 2690 11456
rect 2370 10368 2690 11392
rect 2370 10304 2378 10368
rect 2442 10304 2458 10368
rect 2522 10304 2538 10368
rect 2602 10304 2618 10368
rect 2682 10304 2690 10368
rect 2370 9434 2690 10304
rect 2370 9280 2412 9434
rect 2648 9280 2690 9434
rect 2370 9216 2378 9280
rect 2682 9216 2690 9280
rect 2370 9198 2412 9216
rect 2648 9198 2690 9216
rect 2370 8192 2690 9198
rect 2370 8128 2378 8192
rect 2442 8128 2458 8192
rect 2522 8128 2538 8192
rect 2602 8128 2618 8192
rect 2682 8128 2690 8192
rect 2370 7104 2690 8128
rect 2370 7040 2378 7104
rect 2442 7040 2458 7104
rect 2522 7040 2538 7104
rect 2602 7040 2618 7104
rect 2682 7040 2690 7104
rect 2370 6578 2690 7040
rect 2370 6342 2412 6578
rect 2648 6342 2690 6578
rect 2370 6016 2690 6342
rect 2370 5952 2378 6016
rect 2442 5952 2458 6016
rect 2522 5952 2538 6016
rect 2602 5952 2618 6016
rect 2682 5952 2690 6016
rect 2370 4928 2690 5952
rect 2370 4864 2378 4928
rect 2442 4864 2458 4928
rect 2522 4864 2538 4928
rect 2602 4864 2618 4928
rect 2682 4864 2690 4928
rect 2370 3840 2690 4864
rect 2370 3776 2378 3840
rect 2442 3776 2458 3840
rect 2522 3776 2538 3840
rect 2602 3776 2618 3840
rect 2682 3776 2690 3840
rect 2370 3722 2690 3776
rect 2370 3486 2412 3722
rect 2648 3486 2690 3722
rect 2370 2752 2690 3486
rect 2370 2688 2378 2752
rect 2442 2688 2458 2752
rect 2522 2688 2538 2752
rect 2602 2688 2618 2752
rect 2682 2688 2690 2752
rect 2370 2128 2690 2688
rect 3030 13088 3350 13648
rect 3030 13024 3038 13088
rect 3102 13024 3118 13088
rect 3182 13024 3198 13088
rect 3262 13024 3278 13088
rect 3342 13024 3350 13088
rect 3030 12950 3350 13024
rect 3030 12714 3072 12950
rect 3308 12714 3350 12950
rect 3030 12000 3350 12714
rect 3030 11936 3038 12000
rect 3102 11936 3118 12000
rect 3182 11936 3198 12000
rect 3262 11936 3278 12000
rect 3342 11936 3350 12000
rect 3030 10912 3350 11936
rect 3030 10848 3038 10912
rect 3102 10848 3118 10912
rect 3182 10848 3198 10912
rect 3262 10848 3278 10912
rect 3342 10848 3350 10912
rect 3030 10094 3350 10848
rect 3030 9858 3072 10094
rect 3308 9858 3350 10094
rect 3030 9824 3350 9858
rect 3030 9760 3038 9824
rect 3102 9760 3118 9824
rect 3182 9760 3198 9824
rect 3262 9760 3278 9824
rect 3342 9760 3350 9824
rect 3030 8736 3350 9760
rect 3030 8672 3038 8736
rect 3102 8672 3118 8736
rect 3182 8672 3198 8736
rect 3262 8672 3278 8736
rect 3342 8672 3350 8736
rect 3030 7648 3350 8672
rect 3030 7584 3038 7648
rect 3102 7584 3118 7648
rect 3182 7584 3198 7648
rect 3262 7584 3278 7648
rect 3342 7584 3350 7648
rect 3030 7238 3350 7584
rect 3030 7002 3072 7238
rect 3308 7002 3350 7238
rect 3030 6560 3350 7002
rect 3030 6496 3038 6560
rect 3102 6496 3118 6560
rect 3182 6496 3198 6560
rect 3262 6496 3278 6560
rect 3342 6496 3350 6560
rect 3030 5472 3350 6496
rect 3030 5408 3038 5472
rect 3102 5408 3118 5472
rect 3182 5408 3198 5472
rect 3262 5408 3278 5472
rect 3342 5408 3350 5472
rect 3030 4384 3350 5408
rect 3030 4320 3038 4384
rect 3102 4382 3118 4384
rect 3182 4382 3198 4384
rect 3262 4382 3278 4384
rect 3342 4320 3350 4384
rect 3030 4146 3072 4320
rect 3308 4146 3350 4320
rect 3030 3296 3350 4146
rect 3030 3232 3038 3296
rect 3102 3232 3118 3296
rect 3182 3232 3198 3296
rect 3262 3232 3278 3296
rect 3342 3232 3350 3296
rect 3030 2208 3350 3232
rect 3030 2144 3038 2208
rect 3102 2144 3118 2208
rect 3182 2144 3198 2208
rect 3262 2144 3278 2208
rect 3342 2144 3350 2208
rect 3030 2128 3350 2144
rect 5222 13632 5542 13648
rect 5222 13568 5230 13632
rect 5294 13568 5310 13632
rect 5374 13568 5390 13632
rect 5454 13568 5470 13632
rect 5534 13568 5542 13632
rect 5222 12544 5542 13568
rect 5222 12480 5230 12544
rect 5294 12480 5310 12544
rect 5374 12480 5390 12544
rect 5454 12480 5470 12544
rect 5534 12480 5542 12544
rect 5222 12290 5542 12480
rect 5222 12054 5264 12290
rect 5500 12054 5542 12290
rect 5222 11456 5542 12054
rect 5222 11392 5230 11456
rect 5294 11392 5310 11456
rect 5374 11392 5390 11456
rect 5454 11392 5470 11456
rect 5534 11392 5542 11456
rect 5222 10368 5542 11392
rect 5222 10304 5230 10368
rect 5294 10304 5310 10368
rect 5374 10304 5390 10368
rect 5454 10304 5470 10368
rect 5534 10304 5542 10368
rect 5222 9434 5542 10304
rect 5222 9280 5264 9434
rect 5500 9280 5542 9434
rect 5222 9216 5230 9280
rect 5534 9216 5542 9280
rect 5222 9198 5264 9216
rect 5500 9198 5542 9216
rect 5222 8192 5542 9198
rect 5222 8128 5230 8192
rect 5294 8128 5310 8192
rect 5374 8128 5390 8192
rect 5454 8128 5470 8192
rect 5534 8128 5542 8192
rect 5222 7104 5542 8128
rect 5222 7040 5230 7104
rect 5294 7040 5310 7104
rect 5374 7040 5390 7104
rect 5454 7040 5470 7104
rect 5534 7040 5542 7104
rect 5222 6578 5542 7040
rect 5222 6342 5264 6578
rect 5500 6342 5542 6578
rect 5222 6016 5542 6342
rect 5222 5952 5230 6016
rect 5294 5952 5310 6016
rect 5374 5952 5390 6016
rect 5454 5952 5470 6016
rect 5534 5952 5542 6016
rect 5222 4928 5542 5952
rect 5222 4864 5230 4928
rect 5294 4864 5310 4928
rect 5374 4864 5390 4928
rect 5454 4864 5470 4928
rect 5534 4864 5542 4928
rect 5222 3840 5542 4864
rect 5222 3776 5230 3840
rect 5294 3776 5310 3840
rect 5374 3776 5390 3840
rect 5454 3776 5470 3840
rect 5534 3776 5542 3840
rect 5222 3722 5542 3776
rect 5222 3486 5264 3722
rect 5500 3486 5542 3722
rect 5222 2752 5542 3486
rect 5222 2688 5230 2752
rect 5294 2688 5310 2752
rect 5374 2688 5390 2752
rect 5454 2688 5470 2752
rect 5534 2688 5542 2752
rect 5222 2128 5542 2688
rect 5882 13088 6202 13648
rect 5882 13024 5890 13088
rect 5954 13024 5970 13088
rect 6034 13024 6050 13088
rect 6114 13024 6130 13088
rect 6194 13024 6202 13088
rect 5882 12950 6202 13024
rect 5882 12714 5924 12950
rect 6160 12714 6202 12950
rect 5882 12000 6202 12714
rect 5882 11936 5890 12000
rect 5954 11936 5970 12000
rect 6034 11936 6050 12000
rect 6114 11936 6130 12000
rect 6194 11936 6202 12000
rect 5882 10912 6202 11936
rect 5882 10848 5890 10912
rect 5954 10848 5970 10912
rect 6034 10848 6050 10912
rect 6114 10848 6130 10912
rect 6194 10848 6202 10912
rect 5882 10094 6202 10848
rect 5882 9858 5924 10094
rect 6160 9858 6202 10094
rect 5882 9824 6202 9858
rect 5882 9760 5890 9824
rect 5954 9760 5970 9824
rect 6034 9760 6050 9824
rect 6114 9760 6130 9824
rect 6194 9760 6202 9824
rect 5882 8736 6202 9760
rect 5882 8672 5890 8736
rect 5954 8672 5970 8736
rect 6034 8672 6050 8736
rect 6114 8672 6130 8736
rect 6194 8672 6202 8736
rect 5882 7648 6202 8672
rect 5882 7584 5890 7648
rect 5954 7584 5970 7648
rect 6034 7584 6050 7648
rect 6114 7584 6130 7648
rect 6194 7584 6202 7648
rect 5882 7238 6202 7584
rect 5882 7002 5924 7238
rect 6160 7002 6202 7238
rect 5882 6560 6202 7002
rect 5882 6496 5890 6560
rect 5954 6496 5970 6560
rect 6034 6496 6050 6560
rect 6114 6496 6130 6560
rect 6194 6496 6202 6560
rect 5882 5472 6202 6496
rect 5882 5408 5890 5472
rect 5954 5408 5970 5472
rect 6034 5408 6050 5472
rect 6114 5408 6130 5472
rect 6194 5408 6202 5472
rect 5882 4384 6202 5408
rect 5882 4320 5890 4384
rect 5954 4382 5970 4384
rect 6034 4382 6050 4384
rect 6114 4382 6130 4384
rect 6194 4320 6202 4384
rect 5882 4146 5924 4320
rect 6160 4146 6202 4320
rect 5882 3296 6202 4146
rect 5882 3232 5890 3296
rect 5954 3232 5970 3296
rect 6034 3232 6050 3296
rect 6114 3232 6130 3296
rect 6194 3232 6202 3296
rect 5882 2208 6202 3232
rect 5882 2144 5890 2208
rect 5954 2144 5970 2208
rect 6034 2144 6050 2208
rect 6114 2144 6130 2208
rect 6194 2144 6202 2208
rect 5882 2128 6202 2144
rect 8074 13632 8394 13648
rect 8074 13568 8082 13632
rect 8146 13568 8162 13632
rect 8226 13568 8242 13632
rect 8306 13568 8322 13632
rect 8386 13568 8394 13632
rect 8074 12544 8394 13568
rect 8074 12480 8082 12544
rect 8146 12480 8162 12544
rect 8226 12480 8242 12544
rect 8306 12480 8322 12544
rect 8386 12480 8394 12544
rect 8074 12290 8394 12480
rect 8074 12054 8116 12290
rect 8352 12054 8394 12290
rect 8074 11456 8394 12054
rect 8074 11392 8082 11456
rect 8146 11392 8162 11456
rect 8226 11392 8242 11456
rect 8306 11392 8322 11456
rect 8386 11392 8394 11456
rect 8074 10368 8394 11392
rect 8074 10304 8082 10368
rect 8146 10304 8162 10368
rect 8226 10304 8242 10368
rect 8306 10304 8322 10368
rect 8386 10304 8394 10368
rect 8074 9434 8394 10304
rect 8074 9280 8116 9434
rect 8352 9280 8394 9434
rect 8074 9216 8082 9280
rect 8386 9216 8394 9280
rect 8074 9198 8116 9216
rect 8352 9198 8394 9216
rect 8074 8192 8394 9198
rect 8074 8128 8082 8192
rect 8146 8128 8162 8192
rect 8226 8128 8242 8192
rect 8306 8128 8322 8192
rect 8386 8128 8394 8192
rect 8074 7104 8394 8128
rect 8074 7040 8082 7104
rect 8146 7040 8162 7104
rect 8226 7040 8242 7104
rect 8306 7040 8322 7104
rect 8386 7040 8394 7104
rect 8074 6578 8394 7040
rect 8074 6342 8116 6578
rect 8352 6342 8394 6578
rect 8074 6016 8394 6342
rect 8074 5952 8082 6016
rect 8146 5952 8162 6016
rect 8226 5952 8242 6016
rect 8306 5952 8322 6016
rect 8386 5952 8394 6016
rect 8074 4928 8394 5952
rect 8074 4864 8082 4928
rect 8146 4864 8162 4928
rect 8226 4864 8242 4928
rect 8306 4864 8322 4928
rect 8386 4864 8394 4928
rect 8074 3840 8394 4864
rect 8074 3776 8082 3840
rect 8146 3776 8162 3840
rect 8226 3776 8242 3840
rect 8306 3776 8322 3840
rect 8386 3776 8394 3840
rect 8074 3722 8394 3776
rect 8074 3486 8116 3722
rect 8352 3486 8394 3722
rect 8074 2752 8394 3486
rect 8074 2688 8082 2752
rect 8146 2688 8162 2752
rect 8226 2688 8242 2752
rect 8306 2688 8322 2752
rect 8386 2688 8394 2752
rect 8074 2128 8394 2688
rect 8734 13088 9054 13648
rect 8734 13024 8742 13088
rect 8806 13024 8822 13088
rect 8886 13024 8902 13088
rect 8966 13024 8982 13088
rect 9046 13024 9054 13088
rect 8734 12950 9054 13024
rect 8734 12714 8776 12950
rect 9012 12714 9054 12950
rect 8734 12000 9054 12714
rect 8734 11936 8742 12000
rect 8806 11936 8822 12000
rect 8886 11936 8902 12000
rect 8966 11936 8982 12000
rect 9046 11936 9054 12000
rect 8734 10912 9054 11936
rect 8734 10848 8742 10912
rect 8806 10848 8822 10912
rect 8886 10848 8902 10912
rect 8966 10848 8982 10912
rect 9046 10848 9054 10912
rect 8734 10094 9054 10848
rect 8734 9858 8776 10094
rect 9012 9858 9054 10094
rect 8734 9824 9054 9858
rect 8734 9760 8742 9824
rect 8806 9760 8822 9824
rect 8886 9760 8902 9824
rect 8966 9760 8982 9824
rect 9046 9760 9054 9824
rect 8734 8736 9054 9760
rect 8734 8672 8742 8736
rect 8806 8672 8822 8736
rect 8886 8672 8902 8736
rect 8966 8672 8982 8736
rect 9046 8672 9054 8736
rect 8734 7648 9054 8672
rect 8734 7584 8742 7648
rect 8806 7584 8822 7648
rect 8886 7584 8902 7648
rect 8966 7584 8982 7648
rect 9046 7584 9054 7648
rect 8734 7238 9054 7584
rect 8734 7002 8776 7238
rect 9012 7002 9054 7238
rect 8734 6560 9054 7002
rect 8734 6496 8742 6560
rect 8806 6496 8822 6560
rect 8886 6496 8902 6560
rect 8966 6496 8982 6560
rect 9046 6496 9054 6560
rect 8734 5472 9054 6496
rect 8734 5408 8742 5472
rect 8806 5408 8822 5472
rect 8886 5408 8902 5472
rect 8966 5408 8982 5472
rect 9046 5408 9054 5472
rect 8734 4384 9054 5408
rect 8734 4320 8742 4384
rect 8806 4382 8822 4384
rect 8886 4382 8902 4384
rect 8966 4382 8982 4384
rect 9046 4320 9054 4384
rect 8734 4146 8776 4320
rect 9012 4146 9054 4320
rect 8734 3296 9054 4146
rect 8734 3232 8742 3296
rect 8806 3232 8822 3296
rect 8886 3232 8902 3296
rect 8966 3232 8982 3296
rect 9046 3232 9054 3296
rect 8734 2208 9054 3232
rect 8734 2144 8742 2208
rect 8806 2144 8822 2208
rect 8886 2144 8902 2208
rect 8966 2144 8982 2208
rect 9046 2144 9054 2208
rect 8734 2128 9054 2144
rect 10926 13632 11246 13648
rect 10926 13568 10934 13632
rect 10998 13568 11014 13632
rect 11078 13568 11094 13632
rect 11158 13568 11174 13632
rect 11238 13568 11246 13632
rect 10926 12544 11246 13568
rect 10926 12480 10934 12544
rect 10998 12480 11014 12544
rect 11078 12480 11094 12544
rect 11158 12480 11174 12544
rect 11238 12480 11246 12544
rect 10926 12290 11246 12480
rect 10926 12054 10968 12290
rect 11204 12054 11246 12290
rect 10926 11456 11246 12054
rect 10926 11392 10934 11456
rect 10998 11392 11014 11456
rect 11078 11392 11094 11456
rect 11158 11392 11174 11456
rect 11238 11392 11246 11456
rect 10926 10368 11246 11392
rect 10926 10304 10934 10368
rect 10998 10304 11014 10368
rect 11078 10304 11094 10368
rect 11158 10304 11174 10368
rect 11238 10304 11246 10368
rect 10926 9434 11246 10304
rect 10926 9280 10968 9434
rect 11204 9280 11246 9434
rect 10926 9216 10934 9280
rect 11238 9216 11246 9280
rect 10926 9198 10968 9216
rect 11204 9198 11246 9216
rect 10926 8192 11246 9198
rect 10926 8128 10934 8192
rect 10998 8128 11014 8192
rect 11078 8128 11094 8192
rect 11158 8128 11174 8192
rect 11238 8128 11246 8192
rect 10926 7104 11246 8128
rect 10926 7040 10934 7104
rect 10998 7040 11014 7104
rect 11078 7040 11094 7104
rect 11158 7040 11174 7104
rect 11238 7040 11246 7104
rect 10926 6578 11246 7040
rect 10926 6342 10968 6578
rect 11204 6342 11246 6578
rect 10926 6016 11246 6342
rect 10926 5952 10934 6016
rect 10998 5952 11014 6016
rect 11078 5952 11094 6016
rect 11158 5952 11174 6016
rect 11238 5952 11246 6016
rect 10926 4928 11246 5952
rect 10926 4864 10934 4928
rect 10998 4864 11014 4928
rect 11078 4864 11094 4928
rect 11158 4864 11174 4928
rect 11238 4864 11246 4928
rect 10926 3840 11246 4864
rect 10926 3776 10934 3840
rect 10998 3776 11014 3840
rect 11078 3776 11094 3840
rect 11158 3776 11174 3840
rect 11238 3776 11246 3840
rect 10926 3722 11246 3776
rect 10926 3486 10968 3722
rect 11204 3486 11246 3722
rect 10926 2752 11246 3486
rect 10926 2688 10934 2752
rect 10998 2688 11014 2752
rect 11078 2688 11094 2752
rect 11158 2688 11174 2752
rect 11238 2688 11246 2752
rect 10926 2128 11246 2688
rect 11586 13088 11906 13648
rect 11586 13024 11594 13088
rect 11658 13024 11674 13088
rect 11738 13024 11754 13088
rect 11818 13024 11834 13088
rect 11898 13024 11906 13088
rect 11586 12950 11906 13024
rect 11586 12714 11628 12950
rect 11864 12714 11906 12950
rect 11586 12000 11906 12714
rect 11586 11936 11594 12000
rect 11658 11936 11674 12000
rect 11738 11936 11754 12000
rect 11818 11936 11834 12000
rect 11898 11936 11906 12000
rect 11586 10912 11906 11936
rect 11586 10848 11594 10912
rect 11658 10848 11674 10912
rect 11738 10848 11754 10912
rect 11818 10848 11834 10912
rect 11898 10848 11906 10912
rect 11586 10094 11906 10848
rect 11586 9858 11628 10094
rect 11864 9858 11906 10094
rect 11586 9824 11906 9858
rect 11586 9760 11594 9824
rect 11658 9760 11674 9824
rect 11738 9760 11754 9824
rect 11818 9760 11834 9824
rect 11898 9760 11906 9824
rect 11586 8736 11906 9760
rect 11586 8672 11594 8736
rect 11658 8672 11674 8736
rect 11738 8672 11754 8736
rect 11818 8672 11834 8736
rect 11898 8672 11906 8736
rect 11586 7648 11906 8672
rect 11586 7584 11594 7648
rect 11658 7584 11674 7648
rect 11738 7584 11754 7648
rect 11818 7584 11834 7648
rect 11898 7584 11906 7648
rect 11586 7238 11906 7584
rect 11586 7002 11628 7238
rect 11864 7002 11906 7238
rect 11586 6560 11906 7002
rect 11586 6496 11594 6560
rect 11658 6496 11674 6560
rect 11738 6496 11754 6560
rect 11818 6496 11834 6560
rect 11898 6496 11906 6560
rect 11586 5472 11906 6496
rect 11586 5408 11594 5472
rect 11658 5408 11674 5472
rect 11738 5408 11754 5472
rect 11818 5408 11834 5472
rect 11898 5408 11906 5472
rect 11586 4384 11906 5408
rect 11586 4320 11594 4384
rect 11658 4382 11674 4384
rect 11738 4382 11754 4384
rect 11818 4382 11834 4384
rect 11898 4320 11906 4384
rect 11586 4146 11628 4320
rect 11864 4146 11906 4320
rect 11586 3296 11906 4146
rect 11586 3232 11594 3296
rect 11658 3232 11674 3296
rect 11738 3232 11754 3296
rect 11818 3232 11834 3296
rect 11898 3232 11906 3296
rect 11586 2208 11906 3232
rect 11586 2144 11594 2208
rect 11658 2144 11674 2208
rect 11738 2144 11754 2208
rect 11818 2144 11834 2208
rect 11898 2144 11906 2208
rect 11586 2128 11906 2144
<< via4 >>
rect 2412 12054 2648 12290
rect 2412 9280 2648 9434
rect 2412 9216 2442 9280
rect 2442 9216 2458 9280
rect 2458 9216 2522 9280
rect 2522 9216 2538 9280
rect 2538 9216 2602 9280
rect 2602 9216 2618 9280
rect 2618 9216 2648 9280
rect 2412 9198 2648 9216
rect 2412 6342 2648 6578
rect 2412 3486 2648 3722
rect 3072 12714 3308 12950
rect 3072 9858 3308 10094
rect 3072 7002 3308 7238
rect 3072 4320 3102 4382
rect 3102 4320 3118 4382
rect 3118 4320 3182 4382
rect 3182 4320 3198 4382
rect 3198 4320 3262 4382
rect 3262 4320 3278 4382
rect 3278 4320 3308 4382
rect 3072 4146 3308 4320
rect 5264 12054 5500 12290
rect 5264 9280 5500 9434
rect 5264 9216 5294 9280
rect 5294 9216 5310 9280
rect 5310 9216 5374 9280
rect 5374 9216 5390 9280
rect 5390 9216 5454 9280
rect 5454 9216 5470 9280
rect 5470 9216 5500 9280
rect 5264 9198 5500 9216
rect 5264 6342 5500 6578
rect 5264 3486 5500 3722
rect 5924 12714 6160 12950
rect 5924 9858 6160 10094
rect 5924 7002 6160 7238
rect 5924 4320 5954 4382
rect 5954 4320 5970 4382
rect 5970 4320 6034 4382
rect 6034 4320 6050 4382
rect 6050 4320 6114 4382
rect 6114 4320 6130 4382
rect 6130 4320 6160 4382
rect 5924 4146 6160 4320
rect 8116 12054 8352 12290
rect 8116 9280 8352 9434
rect 8116 9216 8146 9280
rect 8146 9216 8162 9280
rect 8162 9216 8226 9280
rect 8226 9216 8242 9280
rect 8242 9216 8306 9280
rect 8306 9216 8322 9280
rect 8322 9216 8352 9280
rect 8116 9198 8352 9216
rect 8116 6342 8352 6578
rect 8116 3486 8352 3722
rect 8776 12714 9012 12950
rect 8776 9858 9012 10094
rect 8776 7002 9012 7238
rect 8776 4320 8806 4382
rect 8806 4320 8822 4382
rect 8822 4320 8886 4382
rect 8886 4320 8902 4382
rect 8902 4320 8966 4382
rect 8966 4320 8982 4382
rect 8982 4320 9012 4382
rect 8776 4146 9012 4320
rect 10968 12054 11204 12290
rect 10968 9280 11204 9434
rect 10968 9216 10998 9280
rect 10998 9216 11014 9280
rect 11014 9216 11078 9280
rect 11078 9216 11094 9280
rect 11094 9216 11158 9280
rect 11158 9216 11174 9280
rect 11174 9216 11204 9280
rect 10968 9198 11204 9216
rect 10968 6342 11204 6578
rect 10968 3486 11204 3722
rect 11628 12714 11864 12950
rect 11628 9858 11864 10094
rect 11628 7002 11864 7238
rect 11628 4320 11658 4382
rect 11658 4320 11674 4382
rect 11674 4320 11738 4382
rect 11738 4320 11754 4382
rect 11754 4320 11818 4382
rect 11818 4320 11834 4382
rect 11834 4320 11864 4382
rect 11628 4146 11864 4320
<< metal5 >>
rect 1056 12950 12560 12992
rect 1056 12714 3072 12950
rect 3308 12714 5924 12950
rect 6160 12714 8776 12950
rect 9012 12714 11628 12950
rect 11864 12714 12560 12950
rect 1056 12672 12560 12714
rect 1056 12290 12560 12332
rect 1056 12054 2412 12290
rect 2648 12054 5264 12290
rect 5500 12054 8116 12290
rect 8352 12054 10968 12290
rect 11204 12054 12560 12290
rect 1056 12012 12560 12054
rect 1056 10094 12560 10136
rect 1056 9858 3072 10094
rect 3308 9858 5924 10094
rect 6160 9858 8776 10094
rect 9012 9858 11628 10094
rect 11864 9858 12560 10094
rect 1056 9816 12560 9858
rect 1056 9434 12560 9476
rect 1056 9198 2412 9434
rect 2648 9198 5264 9434
rect 5500 9198 8116 9434
rect 8352 9198 10968 9434
rect 11204 9198 12560 9434
rect 1056 9156 12560 9198
rect 1056 7238 12560 7280
rect 1056 7002 3072 7238
rect 3308 7002 5924 7238
rect 6160 7002 8776 7238
rect 9012 7002 11628 7238
rect 11864 7002 12560 7238
rect 1056 6960 12560 7002
rect 1056 6578 12560 6620
rect 1056 6342 2412 6578
rect 2648 6342 5264 6578
rect 5500 6342 8116 6578
rect 8352 6342 10968 6578
rect 11204 6342 12560 6578
rect 1056 6300 12560 6342
rect 1056 4382 12560 4424
rect 1056 4146 3072 4382
rect 3308 4146 5924 4382
rect 6160 4146 8776 4382
rect 9012 4146 11628 4382
rect 11864 4146 12560 4382
rect 1056 4104 12560 4146
rect 1056 3722 12560 3764
rect 1056 3486 2412 3722
rect 2648 3486 5264 3722
rect 5500 3486 8116 3722
rect 8352 3486 10968 3722
rect 11204 3486 12560 3722
rect 1056 3444 12560 3486
use sky130_fd_sc_hd__clkbuf_2  _170_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6532 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2024 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _172_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3680 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _173_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5152 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _174_
timestamp 1704896540
transform 1 0 4876 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _175_
timestamp 1704896540
transform 1 0 7176 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_4  _176_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4232 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  _177_
timestamp 1704896540
transform 1 0 4968 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _178_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _179_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7360 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _180_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9292 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _181_
timestamp 1704896540
transform 1 0 3772 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _182_
timestamp 1704896540
transform 1 0 5428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _183_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1656 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _184_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2668 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _185_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3496 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _187_
timestamp 1704896540
transform -1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2668 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _190_
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _191_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9752 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _192_
timestamp 1704896540
transform -1 0 7176 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7176 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _194_
timestamp 1704896540
transform 1 0 10212 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _195_
timestamp 1704896540
transform 1 0 10304 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _196_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11408 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _197_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _198_
timestamp 1704896540
transform -1 0 3128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2944 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _200_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11408 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _201_
timestamp 1704896540
transform 1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _202_
timestamp 1704896540
transform -1 0 3496 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _203_
timestamp 1704896540
transform -1 0 4784 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _204_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4416 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _205_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3772 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _206_
timestamp 1704896540
transform 1 0 2208 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _207_
timestamp 1704896540
transform 1 0 2576 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _208_
timestamp 1704896540
transform 1 0 3312 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _209_
timestamp 1704896540
transform 1 0 8004 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _210_
timestamp 1704896540
transform 1 0 6992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _211_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3588 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _212_
timestamp 1704896540
transform 1 0 4600 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _213_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _214_
timestamp 1704896540
transform 1 0 4600 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _215_
timestamp 1704896540
transform -1 0 5520 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _216_
timestamp 1704896540
transform 1 0 4508 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _217_
timestamp 1704896540
transform 1 0 5244 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _218_
timestamp 1704896540
transform 1 0 6624 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _219_
timestamp 1704896540
transform 1 0 10120 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 1704896540
transform 1 0 2484 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _221_
timestamp 1704896540
transform -1 0 4140 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _222_
timestamp 1704896540
transform 1 0 10764 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_2  _223_
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _224_
timestamp 1704896540
transform 1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _225_
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _226_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4232 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _227_
timestamp 1704896540
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _228_
timestamp 1704896540
transform -1 0 8372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _229_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _230_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _232_
timestamp 1704896540
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _233_
timestamp 1704896540
transform -1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _234_
timestamp 1704896540
transform 1 0 7728 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _236_
timestamp 1704896540
transform 1 0 6256 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _237_
timestamp 1704896540
transform 1 0 7268 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _238_
timestamp 1704896540
transform 1 0 4876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _239_
timestamp 1704896540
transform 1 0 7636 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _240_
timestamp 1704896540
transform 1 0 8832 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _241_
timestamp 1704896540
transform 1 0 5520 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6992 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _243_
timestamp 1704896540
transform 1 0 10120 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _244_
timestamp 1704896540
transform 1 0 10764 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _245_
timestamp 1704896540
transform -1 0 8464 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _246_
timestamp 1704896540
transform 1 0 8096 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _247_
timestamp 1704896540
transform 1 0 9844 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _249_
timestamp 1704896540
transform 1 0 11040 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _250_
timestamp 1704896540
transform -1 0 11868 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _251_
timestamp 1704896540
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _252_
timestamp 1704896540
transform -1 0 10028 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_4  _253_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10028 0 1 6528
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _254_
timestamp 1704896540
transform -1 0 12052 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _255_
timestamp 1704896540
transform -1 0 8556 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _256_
timestamp 1704896540
transform 1 0 8740 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _257_
timestamp 1704896540
transform -1 0 8740 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _258_
timestamp 1704896540
transform -1 0 11408 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _259_
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _260_
timestamp 1704896540
transform -1 0 10856 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o41a_1  _261_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7084 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _262_
timestamp 1704896540
transform 1 0 7912 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_2  _263_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9752 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1704896540
transform 1 0 10948 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _265_
timestamp 1704896540
transform 1 0 9200 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _266_
timestamp 1704896540
transform 1 0 10672 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _267_
timestamp 1704896540
transform 1 0 10856 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _268_
timestamp 1704896540
transform -1 0 11316 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _269_
timestamp 1704896540
transform -1 0 11960 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _270_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _271_
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _273_
timestamp 1704896540
transform -1 0 8648 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _274_
timestamp 1704896540
transform 1 0 8096 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _275_
timestamp 1704896540
transform 1 0 9476 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _276_
timestamp 1704896540
transform 1 0 9108 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _277_
timestamp 1704896540
transform -1 0 10488 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _278_
timestamp 1704896540
transform 1 0 10764 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _279_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11592 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _280_
timestamp 1704896540
transform 1 0 10396 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _281_
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _282_
timestamp 1704896540
transform 1 0 8188 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _283_
timestamp 1704896540
transform -1 0 8832 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11040 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _285_
timestamp 1704896540
transform 1 0 10120 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _286_
timestamp 1704896540
transform 1 0 7268 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _287_
timestamp 1704896540
transform 1 0 6808 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _288_
timestamp 1704896540
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _289_
timestamp 1704896540
transform 1 0 7728 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_4  _290_
timestamp 1704896540
transform 1 0 8188 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _291_
timestamp 1704896540
transform 1 0 10028 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _292_
timestamp 1704896540
transform -1 0 9936 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o311ai_4  _293_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 11684 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__and3_1  _294_
timestamp 1704896540
transform -1 0 9476 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _295_
timestamp 1704896540
transform 1 0 7360 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _296_
timestamp 1704896540
transform -1 0 7176 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6624 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _298_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9476 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _299_
timestamp 1704896540
transform 1 0 6532 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _300_
timestamp 1704896540
transform -1 0 8188 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _301_
timestamp 1704896540
transform 1 0 7176 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _302_
timestamp 1704896540
transform 1 0 7176 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _303_
timestamp 1704896540
transform -1 0 7820 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _304_
timestamp 1704896540
transform -1 0 8280 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _305_
timestamp 1704896540
transform 1 0 6348 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _306_
timestamp 1704896540
transform 1 0 4692 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _307_
timestamp 1704896540
transform 1 0 5152 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _308_
timestamp 1704896540
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _309_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6348 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _310_
timestamp 1704896540
transform 1 0 5520 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _311_
timestamp 1704896540
transform -1 0 6256 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _312_
timestamp 1704896540
transform 1 0 7360 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _313_
timestamp 1704896540
transform -1 0 6256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _314_
timestamp 1704896540
transform -1 0 5060 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _315_
timestamp 1704896540
transform 1 0 5796 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _316_
timestamp 1704896540
transform -1 0 5428 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _317_
timestamp 1704896540
transform -1 0 6072 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _318_
timestamp 1704896540
transform 1 0 5060 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _319_
timestamp 1704896540
transform 1 0 3772 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _320_
timestamp 1704896540
transform -1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _321_
timestamp 1704896540
transform -1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _322_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5244 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _323_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5244 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _324_
timestamp 1704896540
transform 1 0 4508 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _325_
timestamp 1704896540
transform 1 0 2300 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _326_
timestamp 1704896540
transform -1 0 3128 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _327_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _328_
timestamp 1704896540
transform 1 0 2576 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _329_
timestamp 1704896540
transform -1 0 2760 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _330_
timestamp 1704896540
transform -1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _331_
timestamp 1704896540
transform 1 0 4140 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _332_
timestamp 1704896540
transform 1 0 1472 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _333_
timestamp 1704896540
transform -1 0 3680 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _334_
timestamp 1704896540
transform 1 0 2116 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _335_
timestamp 1704896540
transform -1 0 2944 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _336_
timestamp 1704896540
transform 1 0 2576 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _337_
timestamp 1704896540
transform 1 0 2760 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _338_
timestamp 1704896540
transform 1 0 2024 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _339_
timestamp 1704896540
transform 1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _340_
timestamp 1704896540
transform 1 0 10396 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _341_
timestamp 1704896540
transform 1 0 9752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _342_
timestamp 1704896540
transform 1 0 3772 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _343_
timestamp 1704896540
transform 1 0 4784 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _344_
timestamp 1704896540
transform -1 0 5520 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _345_
timestamp 1704896540
transform 1 0 5612 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _346_
timestamp 1704896540
transform -1 0 5612 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _347_
timestamp 1704896540
transform -1 0 5888 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _348_
timestamp 1704896540
transform 1 0 4968 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_33
timestamp 1704896540
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_44 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_100
timestamp 1704896540
transform 1 0 10304 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_46
timestamp 1704896540
transform 1 0 5336 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1704896540
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_60
timestamp 1704896540
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_84
timestamp 1704896540
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_91
timestamp 1704896540
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_101
timestamp 1704896540
transform 1 0 10396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_110
timestamp 1704896540
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_63
timestamp 1704896540
transform 1 0 6900 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_73
timestamp 1704896540
transform 1 0 7820 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 1704896540
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_115 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11684 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_36
timestamp 1704896540
transform 1 0 4416 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_78
timestamp 1704896540
transform 1 0 8280 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_90
timestamp 1704896540
transform 1 0 9384 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_96
timestamp 1704896540
transform 1 0 9936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_118
timestamp 1704896540
transform 1 0 11960 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_22
timestamp 1704896540
transform 1 0 3128 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_33
timestamp 1704896540
transform 1 0 4140 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_45
timestamp 1704896540
transform 1 0 5244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_57
timestamp 1704896540
transform 1 0 6348 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_65
timestamp 1704896540
transform 1 0 7084 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_89
timestamp 1704896540
transform 1 0 9292 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_97
timestamp 1704896540
transform 1 0 10028 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_110
timestamp 1704896540
transform 1 0 11224 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_118
timestamp 1704896540
transform 1 0 11960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_7
timestamp 1704896540
transform 1 0 1748 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_48
timestamp 1704896540
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_57
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_73
timestamp 1704896540
transform 1 0 7820 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_84
timestamp 1704896540
transform 1 0 8832 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_96
timestamp 1704896540
transform 1 0 9936 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_108
timestamp 1704896540
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_7
timestamp 1704896540
transform 1 0 1748 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1704896540
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_37
timestamp 1704896540
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_58
timestamp 1704896540
transform 1 0 6440 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_73
timestamp 1704896540
transform 1 0 7820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_81
timestamp 1704896540
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_97
timestamp 1704896540
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_9
timestamp 1704896540
transform 1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_33
timestamp 1704896540
transform 1 0 4140 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1704896540
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_90
timestamp 1704896540
transform 1 0 9384 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_119
timestamp 1704896540
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1704896540
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_48
timestamp 1704896540
transform 1 0 5520 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_60
timestamp 1704896540
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_64
timestamp 1704896540
transform 1 0 6992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_74
timestamp 1704896540
transform 1 0 7912 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_91
timestamp 1704896540
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_10
timestamp 1704896540
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_25
timestamp 1704896540
transform 1 0 3404 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_37
timestamp 1704896540
transform 1 0 4508 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_41
timestamp 1704896540
transform 1 0 4876 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_80
timestamp 1704896540
transform 1 0 8464 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_92
timestamp 1704896540
transform 1 0 9568 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_117
timestamp 1704896540
transform 1 0 11868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_11
timestamp 1704896540
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_20
timestamp 1704896540
transform 1 0 2944 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_48
timestamp 1704896540
transform 1 0 5520 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_60
timestamp 1704896540
transform 1 0 6624 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_75
timestamp 1704896540
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_97
timestamp 1704896540
transform 1 0 10028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_104
timestamp 1704896540
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_117
timestamp 1704896540
transform 1 0 11868 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_26
timestamp 1704896540
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_40
timestamp 1704896540
transform 1 0 4784 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_69
timestamp 1704896540
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_82
timestamp 1704896540
transform 1 0 8648 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_88
timestamp 1704896540
transform 1 0 9200 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_97
timestamp 1704896540
transform 1 0 10028 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_117
timestamp 1704896540
transform 1 0 11868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_35
timestamp 1704896540
transform 1 0 4324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_50
timestamp 1704896540
transform 1 0 5704 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_58
timestamp 1704896540
transform 1 0 6440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_66
timestamp 1704896540
transform 1 0 7176 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_72
timestamp 1704896540
transform 1 0 7728 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 1704896540
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_92
timestamp 1704896540
transform 1 0 9568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_113
timestamp 1704896540
transform 1 0 11500 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_17
timestamp 1704896540
transform 1 0 2668 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_25
timestamp 1704896540
transform 1 0 3404 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_37
timestamp 1704896540
transform 1 0 4508 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_72
timestamp 1704896540
transform 1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_79
timestamp 1704896540
transform 1 0 8372 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_91
timestamp 1704896540
transform 1 0 9476 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_103
timestamp 1704896540
transform 1 0 10580 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1704896540
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_15
timestamp 1704896540
transform 1 0 2484 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1704896540
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_61
timestamp 1704896540
transform 1 0 6716 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_66
timestamp 1704896540
transform 1 0 7176 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_78
timestamp 1704896540
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_97
timestamp 1704896540
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1704896540
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_3
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_11
timestamp 1704896540
transform 1 0 2116 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_20
timestamp 1704896540
transform 1 0 2944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_34
timestamp 1704896540
transform 1 0 4232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_40
timestamp 1704896540
transform 1 0 4784 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_45
timestamp 1704896540
transform 1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_53
timestamp 1704896540
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_63
timestamp 1704896540
transform 1 0 6900 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_70
timestamp 1704896540
transform 1 0 7544 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_82
timestamp 1704896540
transform 1 0 8648 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_94
timestamp 1704896540
transform 1 0 9752 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_103
timestamp 1704896540
transform 1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_6
timestamp 1704896540
transform 1 0 1656 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_14
timestamp 1704896540
transform 1 0 2392 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1704896540
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_36
timestamp 1704896540
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_51
timestamp 1704896540
transform 1 0 5796 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_55
timestamp 1704896540
transform 1 0 6164 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1704896540
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_97
timestamp 1704896540
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_114
timestamp 1704896540
transform 1 0 11592 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_120
timestamp 1704896540
transform 1 0 12144 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_7
timestamp 1704896540
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_19
timestamp 1704896540
transform 1 0 2852 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_32
timestamp 1704896540
transform 1 0 4048 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_43
timestamp 1704896540
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_65
timestamp 1704896540
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_75
timestamp 1704896540
transform 1 0 8004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_83
timestamp 1704896540
transform 1 0 8740 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_102
timestamp 1704896540
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_110
timestamp 1704896540
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_113
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_11
timestamp 1704896540
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1704896540
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_54
timestamp 1704896540
transform 1 0 6072 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_67
timestamp 1704896540
transform 1 0 7268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 1704896540
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_96
timestamp 1704896540
transform 1 0 9936 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_108
timestamp 1704896540
transform 1 0 11040 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_120
timestamp 1704896540
transform 1 0 12144 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_7
timestamp 1704896540
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_19
timestamp 1704896540
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_31
timestamp 1704896540
transform 1 0 3956 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_44
timestamp 1704896540
transform 1 0 5152 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_52
timestamp 1704896540
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_67
timestamp 1704896540
transform 1 0 7268 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_78
timestamp 1704896540
transform 1 0 8280 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_91
timestamp 1704896540
transform 1 0 9476 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_103
timestamp 1704896540
transform 1 0 10580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1704896540
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_37
timestamp 1704896540
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_53
timestamp 1704896540
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_57
timestamp 1704896540
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_62
timestamp 1704896540
transform 1 0 6808 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_69
timestamp 1704896540
transform 1 0 7452 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1704896540
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_109
timestamp 1704896540
transform 1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_113
timestamp 1704896540
transform 1 0 11500 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 6532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12236 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1704896540
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1704896540
transform 1 0 7176 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1704896540
transform 1 0 7820 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1704896540
transform -1 0 12236 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1704896540
transform 1 0 9108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1704896540
transform 1 0 7176 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1704896540
transform -1 0 6256 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input19 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1704896540
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1704896540
transform -1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1704896540
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1704896540
transform 1 0 11868 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1704896540
transform 1 0 11868 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1704896540
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1704896540
transform -1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  output28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_21
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_22
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_23
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_24
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_25
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 12512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_26
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 12512 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_27
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_28
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 12512 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_29
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_30
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_31
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 12512 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_32
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 12512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_33
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_34
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 12512 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_35
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 12512 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_36
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 12512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_37
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 12512 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_38
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_39
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 12512 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_40
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 12512 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_41
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 12512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer1
timestamp 1704896540
transform 1 0 4232 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6716 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3
timestamp 1704896540
transform 1 0 6532 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_43
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_44
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_45
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_46
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_47
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_48
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_49
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_50
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_51
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_52
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_53
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_54
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_55
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_56
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_57
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_58
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_59
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_60
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_61
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_62
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_63
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_64
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_65
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_66
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_67
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_68
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_69
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_70
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_71
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_72
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_73
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_74
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_75
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_76
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_77
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_78
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_79
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_80
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_81
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_82
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_83
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_84
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_85
timestamp 1704896540
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_86
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_87
timestamp 1704896540
transform 1 0 11408 0 1 13056
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 A[0]
port 0 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 A[1]
port 1 nsew signal input
flabel metal2 s 4526 14990 4582 15790 0 FreeSans 224 90 0 0 A[2]
port 2 nsew signal input
flabel metal2 s 6458 14990 6514 15790 0 FreeSans 224 90 0 0 A[3]
port 3 nsew signal input
flabel metal3 s 12846 5448 13646 5568 0 FreeSans 480 0 0 0 A[4]
port 4 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 A[5]
port 5 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 A[6]
port 6 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 A[7]
port 7 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 B[0]
port 8 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 B[1]
port 9 nsew signal input
flabel metal2 s 7102 14990 7158 15790 0 FreeSans 224 90 0 0 B[2]
port 10 nsew signal input
flabel metal2 s 7746 14990 7802 15790 0 FreeSans 224 90 0 0 B[3]
port 11 nsew signal input
flabel metal3 s 12846 6808 13646 6928 0 FreeSans 480 0 0 0 B[4]
port 12 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 B[5]
port 13 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 B[6]
port 14 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 B[7]
port 15 nsew signal input
flabel metal4 s 3030 2128 3350 13648 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 5882 2128 6202 13648 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 8734 2128 9054 13648 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 11586 2128 11906 13648 0 FreeSans 1920 90 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 4104 12560 4424 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 6960 12560 7280 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 9816 12560 10136 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal5 s 1056 12672 12560 12992 0 FreeSans 2560 0 0 0 VGND
port 16 nsew ground bidirectional
flabel metal4 s 2370 2128 2690 13648 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 5222 2128 5542 13648 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 8074 2128 8394 13648 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal4 s 10926 2128 11246 13648 0 FreeSans 1920 90 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 3444 12560 3764 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 6300 12560 6620 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 9156 12560 9476 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal5 s 1056 12012 12560 12332 0 FreeSans 2560 0 0 0 VPWR
port 17 nsew power bidirectional
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 opcode[0]
port 18 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 opcode[1]
port 19 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 opcode[2]
port 20 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 out[0]
port 21 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 out[1]
port 22 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 out[2]
port 23 nsew signal output
flabel metal3 s 12846 8848 13646 8968 0 FreeSans 480 0 0 0 out[3]
port 24 nsew signal output
flabel metal3 s 12846 6128 13646 6248 0 FreeSans 480 0 0 0 out[4]
port 25 nsew signal output
flabel metal3 s 12846 4768 13646 4888 0 FreeSans 480 0 0 0 out[5]
port 26 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 out[6]
port 27 nsew signal output
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 out[7]
port 28 nsew signal output
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 out[8]
port 29 nsew signal output
rlabel metal1 6808 13056 6808 13056 0 VGND
rlabel metal1 6808 13600 6808 13600 0 VPWR
rlabel metal3 1050 12308 1050 12308 0 A[0]
rlabel metal3 866 11628 866 11628 0 A[1]
rlabel metal1 4600 13294 4600 13294 0 A[2]
rlabel metal1 6532 13294 6532 13294 0 A[3]
rlabel metal2 12190 5593 12190 5593 0 A[4]
rlabel metal2 9706 1588 9706 1588 0 A[5]
rlabel metal2 8418 1520 8418 1520 0 A[6]
rlabel metal2 6486 1554 6486 1554 0 A[7]
rlabel metal3 820 7548 820 7548 0 B[0]
rlabel metal3 1050 10948 1050 10948 0 B[1]
rlabel metal1 7176 13294 7176 13294 0 B[2]
rlabel metal1 7820 13362 7820 13362 0 B[3]
rlabel via2 12190 6851 12190 6851 0 B[4]
rlabel metal2 9062 1027 9062 1027 0 B[5]
rlabel metal2 7130 1588 7130 1588 0 B[6]
rlabel metal2 5842 1588 5842 1588 0 B[7]
rlabel metal1 6256 12274 6256 12274 0 _000_
rlabel metal1 8602 12274 8602 12274 0 _001_
rlabel metal1 10948 11118 10948 11118 0 _002_
rlabel metal1 11914 7378 11914 7378 0 _003_
rlabel metal1 8418 6766 8418 6766 0 _004_
rlabel metal1 9798 6324 9798 6324 0 _005_
rlabel metal1 11270 5746 11270 5746 0 _006_
rlabel metal1 11086 5712 11086 5712 0 _007_
rlabel metal1 10580 6834 10580 6834 0 _008_
rlabel metal1 11316 7378 11316 7378 0 _009_
rlabel metal2 9982 6970 9982 6970 0 _010_
rlabel metal2 10994 6528 10994 6528 0 _011_
rlabel metal2 12006 6630 12006 6630 0 _012_
rlabel metal1 10902 6256 10902 6256 0 _013_
rlabel metal2 9062 6086 9062 6086 0 _014_
rlabel metal1 8142 6188 8142 6188 0 _015_
rlabel metal1 11178 6324 11178 6324 0 _016_
rlabel metal1 11454 6426 11454 6426 0 _017_
rlabel metal2 10810 6817 10810 6817 0 _018_
rlabel metal2 7498 5066 7498 5066 0 _019_
rlabel metal1 8878 3570 8878 3570 0 _020_
rlabel metal1 10258 3128 10258 3128 0 _021_
rlabel metal1 10902 2992 10902 2992 0 _022_
rlabel metal2 10442 3842 10442 3842 0 _023_
rlabel metal1 10856 3978 10856 3978 0 _024_
rlabel metal1 11822 4148 11822 4148 0 _025_
rlabel metal1 11500 4114 11500 4114 0 _026_
rlabel metal2 11546 4284 11546 4284 0 _027_
rlabel metal1 9522 12104 9522 12104 0 _028_
rlabel metal1 9568 12410 9568 12410 0 _029_
rlabel metal2 7590 11424 7590 11424 0 _030_
rlabel metal2 8510 11492 8510 11492 0 _031_
rlabel metal1 9384 11798 9384 11798 0 _032_
rlabel metal2 9982 11900 9982 11900 0 _033_
rlabel metal1 9706 11662 9706 11662 0 _034_
rlabel metal2 10626 11322 10626 11322 0 _035_
rlabel metal1 11270 12070 11270 12070 0 _036_
rlabel metal1 11040 11186 11040 11186 0 _037_
rlabel metal2 10718 5678 10718 5678 0 _038_
rlabel metal1 8556 4590 8556 4590 0 _039_
rlabel metal1 8050 4794 8050 4794 0 _040_
rlabel metal1 9660 5338 9660 5338 0 _041_
rlabel metal2 10718 5168 10718 5168 0 _042_
rlabel metal1 7038 3570 7038 3570 0 _043_
rlabel metal1 7498 3060 7498 3060 0 _044_
rlabel metal1 7912 2958 7912 2958 0 _045_
rlabel metal1 8234 3026 8234 3026 0 _046_
rlabel metal2 10166 3230 10166 3230 0 _047_
rlabel metal1 9982 4114 9982 4114 0 _048_
rlabel metal2 9246 3366 9246 3366 0 _049_
rlabel metal1 9284 3162 9284 3162 0 _050_
rlabel metal1 8326 3162 8326 3162 0 _051_
rlabel metal1 7268 10030 7268 10030 0 _052_
rlabel metal1 6992 9554 6992 9554 0 _053_
rlabel metal2 6762 9146 6762 9146 0 _054_
rlabel metal1 6854 9044 6854 9044 0 _055_
rlabel metal2 7590 7344 7590 7344 0 _056_
rlabel metal1 7544 4590 7544 4590 0 _057_
rlabel metal1 7452 4794 7452 4794 0 _058_
rlabel metal1 7268 5338 7268 5338 0 _059_
rlabel metal1 7728 4114 7728 4114 0 _060_
rlabel metal1 5014 2924 5014 2924 0 _061_
rlabel metal1 5198 4046 5198 4046 0 _062_
rlabel metal2 6394 3536 6394 3536 0 _063_
rlabel metal2 6302 3128 6302 3128 0 _064_
rlabel metal2 6026 3808 6026 3808 0 _065_
rlabel metal1 5796 3570 5796 3570 0 _066_
rlabel metal2 5842 4828 5842 4828 0 _067_
rlabel metal1 5934 9452 5934 9452 0 _068_
rlabel metal2 5842 7548 5842 7548 0 _069_
rlabel metal1 6118 5712 6118 5712 0 _070_
rlabel metal1 5796 5882 5796 5882 0 _071_
rlabel metal1 5566 6256 5566 6256 0 _072_
rlabel metal2 5658 5984 5658 5984 0 _073_
rlabel metal1 4554 3502 4554 3502 0 _074_
rlabel metal1 4738 3672 4738 3672 0 _075_
rlabel metal1 5934 3604 5934 3604 0 _076_
rlabel metal1 5060 3706 5060 3706 0 _077_
rlabel metal2 4462 3876 4462 3876 0 _078_
rlabel metal1 2530 6664 2530 6664 0 _079_
rlabel metal2 2806 6732 2806 6732 0 _080_
rlabel metal1 3082 6324 3082 6324 0 _081_
rlabel metal2 2622 6596 2622 6596 0 _082_
rlabel metal2 4462 8262 4462 8262 0 _083_
rlabel metal2 4186 8806 4186 8806 0 _084_
rlabel metal1 2438 8398 2438 8398 0 _085_
rlabel metal1 2346 8908 2346 8908 0 _086_
rlabel metal2 2162 8772 2162 8772 0 _087_
rlabel metal2 2990 10200 2990 10200 0 _088_
rlabel metal1 3358 9554 3358 9554 0 _089_
rlabel metal1 2530 8976 2530 8976 0 _090_
rlabel metal1 2668 9146 2668 9146 0 _091_
rlabel metal2 9798 8636 9798 8636 0 _092_
rlabel metal1 9752 8602 9752 8602 0 _093_
rlabel metal1 4830 9690 4830 9690 0 _094_
rlabel metal1 5382 9520 5382 9520 0 _095_
rlabel metal2 5934 8262 5934 8262 0 _096_
rlabel metal1 5014 8432 5014 8432 0 _097_
rlabel metal1 5658 8262 5658 8262 0 _098_
rlabel metal1 5704 9146 5704 9146 0 _099_
rlabel metal1 10350 7820 10350 7820 0 _100_
rlabel metal1 3450 6324 3450 6324 0 _101_
rlabel via2 4922 8483 4922 8483 0 _102_
rlabel metal1 10304 4454 10304 4454 0 _103_
rlabel metal2 9154 8704 9154 8704 0 _104_
rlabel metal1 5198 8568 5198 8568 0 _105_
rlabel metal1 2254 7854 2254 7854 0 _106_
rlabel metal1 6394 7344 6394 7344 0 _107_
rlabel metal2 6578 7718 6578 7718 0 _108_
rlabel metal2 9522 8262 9522 8262 0 _109_
rlabel metal1 11086 8500 11086 8500 0 _110_
rlabel via2 3174 9571 3174 9571 0 _111_
rlabel metal1 2162 7786 2162 7786 0 _112_
rlabel metal1 3496 8398 3496 8398 0 _113_
rlabel metal1 3496 8466 3496 8466 0 _114_
rlabel via1 2162 9078 2162 9078 0 _115_
rlabel metal2 2162 6970 2162 6970 0 _116_
rlabel metal2 2898 8942 2898 8942 0 _117_
rlabel metal1 2346 9554 2346 9554 0 _118_
rlabel via2 2622 9469 2622 9469 0 _119_
rlabel metal1 9890 8976 9890 8976 0 _120_
rlabel metal1 10166 8466 10166 8466 0 _121_
rlabel metal1 7222 7310 7222 7310 0 _122_
rlabel metal1 10350 7480 10350 7480 0 _123_
rlabel metal1 10994 7786 10994 7786 0 _124_
rlabel metal2 10994 7684 10994 7684 0 _125_
rlabel metal1 11178 8432 11178 8432 0 _126_
rlabel metal2 11546 8704 11546 8704 0 _127_
rlabel metal1 3036 5542 3036 5542 0 _128_
rlabel metal1 2300 8466 2300 8466 0 _129_
rlabel metal2 11362 8772 11362 8772 0 _130_
rlabel metal1 2438 12172 2438 12172 0 _131_
rlabel metal1 3404 11730 3404 11730 0 _132_
rlabel metal1 3128 11730 3128 11730 0 _133_
rlabel metal1 3772 11322 3772 11322 0 _134_
rlabel metal1 2530 12240 2530 12240 0 _135_
rlabel metal1 3496 10574 3496 10574 0 _136_
rlabel metal2 2990 10812 2990 10812 0 _137_
rlabel metal2 4830 10064 4830 10064 0 _138_
rlabel metal1 7222 12172 7222 12172 0 _139_
rlabel metal1 6992 12818 6992 12818 0 _140_
rlabel metal1 5244 12818 5244 12818 0 _141_
rlabel metal1 4922 12240 4922 12240 0 _142_
rlabel metal2 5198 12070 5198 12070 0 _143_
rlabel metal1 5152 11322 5152 11322 0 _144_
rlabel metal1 4922 12410 4922 12410 0 _145_
rlabel metal1 5612 12750 5612 12750 0 _146_
rlabel metal1 6762 12682 6762 12682 0 _147_
rlabel metal1 8694 12614 8694 12614 0 _148_
rlabel metal1 10948 10642 10948 10642 0 _149_
rlabel metal1 4186 5678 4186 5678 0 _150_
rlabel metal1 11638 7514 11638 7514 0 _151_
rlabel metal1 10534 10064 10534 10064 0 _152_
rlabel metal1 3174 6732 3174 6732 0 _153_
rlabel metal2 4002 6562 4002 6562 0 _154_
rlabel metal1 5842 8398 5842 8398 0 _155_
rlabel metal2 4830 4998 4830 4998 0 _156_
rlabel metal1 8602 5610 8602 5610 0 _157_
rlabel metal1 8418 8466 8418 8466 0 _158_
rlabel metal2 8050 8772 8050 8772 0 _159_
rlabel metal1 9384 9146 9384 9146 0 _160_
rlabel metal1 11224 8874 11224 8874 0 _161_
rlabel metal1 11132 8942 11132 8942 0 _162_
rlabel metal1 8878 12410 8878 12410 0 _163_
rlabel metal2 5750 11492 5750 11492 0 _164_
rlabel metal1 6992 11730 6992 11730 0 _165_
rlabel metal1 7774 12818 7774 12818 0 _166_
rlabel metal1 8050 12138 8050 12138 0 _167_
rlabel metal1 8694 12750 8694 12750 0 _168_
rlabel metal1 9890 12682 9890 12682 0 _169_
rlabel metal1 1656 12614 1656 12614 0 net1
rlabel metal2 3818 7922 3818 7922 0 net10
rlabel metal1 7314 13158 7314 13158 0 net11
rlabel metal1 7866 13260 7866 13260 0 net12
rlabel metal2 9246 6426 9246 6426 0 net13
rlabel metal1 9338 4590 9338 4590 0 net14
rlabel metal1 7268 2482 7268 2482 0 net15
rlabel metal1 5842 2482 5842 2482 0 net16
rlabel metal2 2254 5440 2254 5440 0 net17
rlabel metal1 2070 5712 2070 5712 0 net18
rlabel metal1 2622 5644 2622 5644 0 net19
rlabel metal1 4600 12206 4600 12206 0 net2
rlabel metal1 1932 6970 1932 6970 0 net20
rlabel metal2 2070 7956 2070 7956 0 net21
rlabel metal1 1702 7888 1702 7888 0 net22
rlabel metal1 11914 9044 11914 9044 0 net23
rlabel metal1 11914 5236 11914 5236 0 net24
rlabel metal2 10166 4998 10166 4998 0 net25
rlabel metal1 8464 2414 8464 2414 0 net26
rlabel metal1 4738 5610 4738 5610 0 net27
rlabel metal1 4600 3910 4600 3910 0 net28
rlabel metal1 5566 5134 5566 5134 0 net29
rlabel metal1 4738 13158 4738 13158 0 net3
rlabel metal2 7958 7548 7958 7548 0 net30
rlabel metal1 6578 3468 6578 3468 0 net31
rlabel metal1 6532 13158 6532 13158 0 net4
rlabel metal1 10672 6290 10672 6290 0 net5
rlabel metal1 10166 2618 10166 2618 0 net6
rlabel metal1 8234 2618 8234 2618 0 net7
rlabel metal1 5842 2618 5842 2618 0 net8
rlabel metal1 5014 7480 5014 7480 0 net9
rlabel metal3 751 4828 751 4828 0 opcode[0]
rlabel metal3 1096 5508 1096 5508 0 opcode[1]
rlabel metal3 751 6188 751 6188 0 opcode[2]
rlabel metal3 1096 6868 1096 6868 0 out[0]
rlabel metal1 1610 8058 1610 8058 0 out[1]
rlabel metal2 1518 8449 1518 8449 0 out[2]
rlabel metal2 12098 8857 12098 8857 0 out[3]
rlabel metal2 12098 5763 12098 5763 0 out[4]
rlabel metal2 11730 4913 11730 4913 0 out[5]
rlabel metal2 7774 1520 7774 1520 0 out[6]
rlabel metal2 5198 1656 5198 1656 0 out[7]
rlabel metal2 4554 1520 4554 1520 0 out[8]
<< properties >>
string FIXED_BBOX 0 0 13646 15790
<< end >>
